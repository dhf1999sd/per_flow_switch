`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kWm9V5Mvg0pGEImXjnz7gpNYOqrR4sCC6H0xDFTz06gdjd+GQTUPGBELgrdfExOSCnors3JMXPXw
0ECTstxBCQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Fcxb4Ecwx1GRn7EPimAplMJJjm5/mEhngx/XMHk56lWshePCfNsPUQLoD4tlX3WJk3JUL35375XJ
omFuoiA1Mb7fDl0P9S1gzjOTjkc/jpNW844eiAYO68cBV/+Ks78DBBGBPwdvJObBzzkVNwQqRhgZ
2WuKH4p1h5qmvJ42WL0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uPXyrd1cFxPIG76cbtiCWWBDYZO+AvDb6GpIEPieUG4goHUaymihtiPk5GcmAOUqqIUu2ffdCGPl
bHEAWfZ3K5QPSHdrnaO2DDNX2Sr/YfxGUf8h4fQ4+PZiViryo5Bxd+qwadw7qJh5wI/FyOir/zik
USP/3nSGAk+LLWIH0ob8bTNGJMpEAtUfcPAGcbOvgG0kNC6ur2D4smbFZNU3xHRjRe3+Q8fkU3EZ
2fgiA8Rj07NJqm5vrmBllX04z2RTY+TWQhuYK8aL/Q5uLkkTPNiMFnbv13pSf2SapZZn4gNPtLfC
phnRbJM8BOgZX3/0RkZ+rg+4oMq2eNfW43mC3Q==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fxi8k2EoO+KEvv1G5caLKoJea3rwiOc75U3qEUlcDP6caNFwRDPPwOe/bkaUvbBxk+7e5gg8F91K
TXyx+lJgdjapbLFFKrjXYK6CPd5KzD3C3aWZlpWvIYDN1NUAMuvGGJf/iv2VwGYdPal4OeWBg4Dz
fyg7vkm6s6UDAaNcTsY+8oETVsbDWOIM4haH9kNsTh+Y6enWUW7VX+dD8WeU+0sx1ZRxgVhvMATR
4lEJp2Rr6bUrHkI9we9b+1dp+coFEG/o6EUHqcL2yE/4gAA8ZAVKabySEDYb+LM8T/8khT256VFP
Upsb1FjWOvDmhJdPVSwb/zGysBQz2o7FLv+JZw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vHRJG9lNgGUgtOANb2urw8ch6tPEovtogAmnKE9HwnfA2yPSWKeYhSmtzdLQfoRfMhDj/OyN9TNL
1EivC0qCpW0Cx8IbyvABcxqRdwXklaOlboj7s4v2wyHCgJgqG4zTLYVc7MqJaVji6FW103obxWnu
TAuL8sL45/hcbGvNiO+3nGiM75KWWxA8qQKHnfxSTh6YW4+9nGwp+ZLgl/P0vrXTfEVkgiGoFjdX
wmHFmy2kSsTkG34YKyJYn2tl+85xHMPqAizEEGbaUOyQc+QOSjsYXB3VHQlQNN2qkn+a944GlwmZ
ANgphbMp6A+3vNLxAfEyV4H5oQ4lnjzJ4gJrBw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
O4GmhGCjYsUqXFQBHHOq3NSDxr1jcAsW9rSpJrrad3qWqiYS7VdUVZBBLANqKvfHNPimxkc7MUg7
Ml9E0bUt51tkCdtcgUENkAMJ17uRx7YMWjGw6IJHx8KGxQ745lXDw1277/f5xUTJih7DALrlnxQZ
aYEUDiK+UU+unU8Y0nU=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
X1toi5TgJlCoO+ockymOLfXcpspFDqUhanzWdxQJrg3OATFpqeEOogtTCzpFhza2xKcGoYzQ3hA8
4B6VxNA8F4/d3pB+5uHPZZYK2xdKdJWE/lWu7UN7D9xVfP8soVc64fh+YoJeh2IQGaA+XgbJq7/l
6k6YstDr3uB5BDIVVSQxXRl8/+6i79w9ottt8E0USMm1JOs73zR6kMu3ccdEkNrSDNyhpbE/fIdm
z4s8OWs2AmCCobL18sGNtIs0C3Bf1PMht8P50o00WTOx1LbhdkCb655ZLnj/D33bI7XaKgPQNDw1
IUxQptpThWCV3vNsp1jSPmC9WYWHPUQmg6geUg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 170448)
`protect data_block
YQnE2aYZT9dbX249nG1+v4FWRLdouivcLg3VVjd0v0glPVvAQhhcys0KWbCXkJ+SlEfBB73oxGTN
aSqGMk/9XA4E6l8JfEY0rlyit7SuwdrkCCWlfqcvbQEbVR7n18VGWPY/jqfSZJbo/gVn8DnmgNua
8hjsBWaQOILbnTqX0HH804HegJRUuV3OX++Rq230cw317qy8RbKgGQZMCrPS7+ujotat9/tHG1cx
EOL+5Rc2NVdedvKTlZHRzLJrWgrqnKu1zxru8dIBRnoPUN5y3e07bXmZw5PCKIs1A3JzK+Jac6MC
lxjsJHCcT5c4NNY6iQiCbs45FO3WYSbrRB38pCUml/zQ5ZIwcxU0bQYNNi8hUkBmLVzsHuGiCgmG
fDxBnCCV2D8eX/2byVHQ5e+dC/BsGDj6PSfQaQ1ZYbDPHx8xFYr8V9gVbOf681o7pYY+AVzLaEoK
I6IiKDxN8NYcyoPQdOppGxrS9qf1t+WfBnmiE+6ROX781b0eX0Rw4br2QZrLuYd0Vto1FC3nLSah
w3MlbPKHaZyi3NGvQ9VdVWB2HiAtHpjJX22DzgJttu/sf1LmPEVokQtCRJvdVC3xZwAdwvBuBF4m
EM00VJXxZoKJF/LRietDMkrE+ba9wUeoQxeB6tSrFCh/Uu+a+sxJK5uiGM+Huv027qm9Dksv3cff
rjJwJRtcQSHGpEOVnndKY1sDV9coaCsYHcPFenQnAreouw3YIqP1yCKelH6YwrHsEnistIJFas11
wUmIta9ma6XSC0FkVSXf7B9KTj6MJ5bLtKNkyAXkucaSaCG8oRj2gGP2tOfhsSHG/1DPNWDxltp9
KKB5LLAZ2ZvuNvtvQ+j95TLf27KKOM8jF17E88CEBTKdabK1rE5wqsV5FLU8PDmJDf+k/jz6VP7f
giYwLwhiEwLdxNlS6gczwASW9v5FLFBb7J/da7LHU6sNgIuT8t75xX4T8rMIHKfR99prJ59QzF5T
fx/IzB+jELagIURkBrnvQvczeBkKbTK8F+q2LhsDgNG+7L2iChCvuT+U3K4j1Cel6OTZRdTkBUai
MOI0/0l3WaItYLJ84I31Cln1VMloT3dZOVqCDarPiIdm6Rq/C3rG57r6gPd/YszYtqybGS7e/Epk
urlXZ35CDgNIEid3lIhGnpSXFffLE5xW/xBtZyHj3iPy7C+HJ0v8+LJqwg3FcohCZk5frM+i24tF
n0n9HTTc4BLz+dJ8qlXTwi3krzOWkkUsc4DI/Y2cHOX6+kQtfoIk0BQOyvsHiMOWRdAJ0o81aulI
89FuHoqv9bLTmSxxKXFjo16TOZMOktC9JbVwP6MlcqQ2sMnkGwk6DtdlkiEYXGztdmESK0Fsd7Lr
QRz/x3yEcm/W5SJGCumAi/toeUXB2zQmHE6bZlkzzXOwUWckgmBLpmkoJ7Jv7tBCWaLJew0YyHAu
WgzY8ccw9kqQtkzDcVCYoIe1vP1YMT3x0nCPE2eLyQrQfyzxAW1DwtnWX1C6Y0GGzzakQKOjAjD0
h6uynBQpLgl45ZF7a2ezZIURsXULq5JNl2C4aWmey8b+qlyWYtjEHkp3qqgGq18UNYl4ED93BZEw
LMdfCKs8/hbbnRV9V6p4V5VKDNBC7da29aGR66DEkc/E+cLmr+a0G2RlK2ZqQxaXTnoFZ61cZ2r8
sOPS1WtTId85mbmbK0BYReLP/k7LPsizdRIvlMSDYEb5BfQLCPsAHGa+ENrZiMtGyBR02ozzxaZ0
5N93dDPh5JV5KB1+KNRLyuM5dQaHnx6AA9Dv7s5zXFNmdIwmdRXUpyMZFijrEERJN9Hy2fWgO0zx
3e3PNmoz58YRRal1530zepyiH5AHMei++Qz+8HTE+gIt5u86ehCa4C+ekoy/tNL90oshAuUG4LmR
od9JwDNY9rGr2AEnZbd+AkAGHlyfTFeQp7268ao7AiqSbQcgQ5SYeGY3hcDvDFQdS7LTbLoCXvNh
C1wwWx9sS/PMqz0zFuPUJi4ag0knR6VdZMU5SX/6mPIlP5oHDVJ3snZzUD9ks/wPx36EfReCPkwQ
IW6SG3hw2MIBysEnJPO7eyO/pj7kJYFhKkurfLUpf4fxcEivyGAK5tYfUWuBfEEhclWbXAT/Gpfb
r+1MqVn8DqQRiNrDUE3wC0O2YaDS7ZT6+uvkft8We8bGBykCMfHlcAv+Rz+0hiozfhHJy7DVONxL
0nkvU4dR1oXnbUE5s2adytlT6pSCcObW9lxBqmWbuz2bwA8sLt+KC7/XzvWG+uONGON2RBFz2ZN3
OSuqm4N5fdPKX/PgoOZfqnuS6Jj0ggRc/LaAhhOit04qTkgm6eM/AUBxFjHlpMPMmKYeAOBL8om/
c21C3R7QUspj7woCG9DUoYePEgPVJsBF1KBySFxvQ92EMMcprODxfloAG4rII6u3QWyuLI4D3ncy
H/FeRyKYsyHbO0HlDtKNnB9GDi0YeLV9BFrk6GebZggbvBGPWcwVwI1Etfwr5Rmk3euuHckip8/k
F4Lrh5OUi/FFHX1KnDT8Wba1VnZDZEziw9Mr0yW6z4YocN4AZoBrw1YXmj7bYaJdaSokx9asFanJ
t7/2ozkcsE4vMmWZfiykht2bRu01dkZB+YPviIrkB1Yue1OuguwGd+PlyvUhN2JliKcw4PkTrKOi
+EDOn0QfPl/sPwK03yy5suDiasHLp/4vI97dnC50tUxJVAREaEAA5krNGTwJKj3MAu5tdc7+UdOQ
V8il8+pAagKSeWdWDGxEtUuisnwv8Ufn1wTDNsQfVUzoqYdkfSDloy5+TMW3026JyxNir62mCYhh
7S/dkfyb1ig/5ygT4I3zSGkIfhI5RX3OOQdS0DZSmYcAuYwGwGkXbyerVw5IZ42kn7J5IXbZnVUF
DT/yb3uXqrr2DVAuTlO4ilRsdjyLZ8jfuWAEFzlRfSlC1x1S+4DYx/rs0yuYhvRBx4xG83Lr/hlv
L0wff2ltl5/pbD9IHVzXMyZNdACB+lpSrpAWv8zEF0zCdhODY6kHTNK+jePilgApX+RBJ0eZ1q8e
PE7tGPzuP7+IgWdCyXFYi01HDi8NyWcrxZ30dtB9Z7cxU7JD0/8VxqfMxivgCCeuy0SpQN8zdgIr
EFL2ckYJnxDRqvcrqYtJxPccHWfRthNSws9z9rM1e8SH5wgrO/N3jmNGGD0EvGSlgRdPr4WUHjNk
uBv3UedVJ0mNDbLDx1mZ2tvpYucC4XpvSoUP8T0Tacrh7Ip+zL5Lt4foFdLQmLTolo1BG+xUjNxs
gnPNl+kv/2pqOmVJtLABMp6jQKhmO8brHjTaCMVMMcbsqOqizLf83veeRiMGSKk8/9NDlKmvT9EF
InpdNyZjq5LPC5eC/EQKiHsYRvpFwTGKKQosp/15EL+K+cpUAMcqOHis4TWXkw24bfDRWLdF+5lH
EP88ZggpuNCrmJvuOVyMl096dp6kN1R5xlijCztmfJWXl5eUXPxOPFNJHwXA6RCDmML6oMIRlKDJ
JyW1VpZjfHtPrRdTz849ifo4zYWIz0k6AQH6G9pUYCRGQVlUSn07fgxZrZX4QZPBfpaxudpb9YN/
+37PyIeB/rI4DYgyBcrh2jlsAuk283UZYcX+1kysB6KTe3RzRlnZxZIiMZVkPZAyk0819N23anFn
v9UvKBZb0gjdHiYLvAFAwsQgSBID1S9ODa/qt9GaDE2t0oEqRP5zRK0Vx66RSfVD72Ucj91aELxk
tzMMwzuKwFmgEoRYQfK4r57/VxDk9EuD6FsnY4T2hOPD+DAbRrW3QeBEkFMk4fTAubRgECRA3rPe
eTnPKn1vg7+8PgUKaeap5Ztm0y8ZDZKcJ9HnczAlFZAzy7iuJ92tV2YSA9B0LctSWvYJme3NN83+
401UzmF8UsCzLMov1ggxmjeH0ZsCpmc9uyy9M9JMusmM/oIizcFN7QwtuMUndpv5EVBulWKrbrLi
sGEBDdnqBeZ6VV46BB+WifvwrP1ZAfEfZW4NQF/uQh24q+hnEimnT61uiaehPWwOsEzdbAKs2njD
Su2QWWkKTFXPxC7Oj4WTsaseogJBeZ1LaHVdc/xjTyuWXjhIhuyWonztNIROZsA7D+pAh7f+2aN1
NrN3Sk9FDw2xXMpXYeHYTYGxjsVQ/08OYkQ6bXBaHPaCBKb39AgY7zdwTTESK961s6ILnizpPabV
uvBU1mPGTDVuGO0RcEcWYeScJwg9GQoTVsSrfnwIUTNVOL8icf3xpdBO41uPU1ZuZzTMbOcfggG4
94BYtIRRrm1anLT+mD/4EbTlWcZClgDTmhBkrWuT0rNg30Ed1abifhk68ewoHFr4dkZmB0Cc5/ga
iCKtp6SfyElNGLQaCRMxEhjZstHbny0Xyak5gowBb1Dks0Gz2gwUy0qyd9Fm5gPubrE3Zoje0Emi
GumUWeq4YFP0d2jlxi3kzDVVmeZz/AJ7NjtUcXcSlfw3RfSV33Ug4MrYk63nu5khv8stWrEgHtg5
pJv+nrfbhHa9N+rmEYSfeBfLP7cgOVvq4j8BT98/NK4qj83kCB267z8j8VDWcEexxTKqXog7Z2he
4301woJvJY9QS9fEtH8eU7adLiNimDKUIvphtF7Nd5eOISR1n3Kuu77hcG12CzRgc1mG1X/0NEvr
L2+3cWO4336G3q9du+qGLqHdoxMAFkVtaN0hqoIW8vC10H5kVBfQX1fJwclPP+0WBOWpF8wq+WlI
41iZ3/rTP/oArcO6Gi8eIY33p/TGcFHG/1nC9BUrt+2AAkCRwBoj/duhy5L3Mh1DCh8wtz8vsXqi
1apRe+05pBiXYWlAkgivdRUu3765y+YzbbEiaH0ISEnskk32twSkRtb7esPkeXLzktPoQRqaefjj
fdNAr+sSOP+pOhJdRFWjeBxiPFvkHhTkkyzbmO06phTtBGGZA0ScroNOkgTnG5a4QKbP2IKnhhDf
kE90N1gRE7H0XUfBaQbOEQbhwqZa/og7mldVwsfC95rrOM5iyLmyU5tZ9r7UV7s5+EzMp0f7CEdQ
lTxck7bfYmJkBmNxNPas2MooJ6cK09st6tltjUD9/4vQjgucSlm99L9QUybH8RwPihoVrBR9XoQc
FF4NqQdJkFFQBPUcBHcMsA+wZ9JH4SpYvpUUkcpFvyESbkkrqtSAEqIcEr1RTYY3HU6avE6Uve+e
iFfIduR/F2/Z8tETaoANABexNfmGh+Gdvie4xnC+STeU4uFoGjsJfPG4wAchABioPQWNl8qFx5Nx
m4oHsKLa9yhLBxEoQvhzoN9j+M0Q8clbFrJsYGNdtOjYpflko/yiV6LIbg1bOORllObGuZ/LW7vT
xa+cKX0XTeHHetMnqiHFkkMk6/ZJ+A2/S9RaEukzyoxoZt5tF+R/svInzN2pTMq8PLAhyTvlEdEV
qYRKcqPxxzNV4vliRhl7TC45ko1dE7I99lJU9AFb/+RzxwJrUs/DDb85sfP8DnpYGUQU2jkBXwn9
4R6PZpvhpuKmvrCnlzT+1kqy4Xq9H9U2e+SHiIEUuX+Hwr2YgPdPzFyCnfz7ip+09rfrkWtORliV
mVkFO/b+64J/+X4Bz95wWdyfH2F+M4Ut7siUKxBNXyKwFSJa0Yu98EDtl0ygN/ogryqML1ZJWLc2
9ost4Trjxjdk8IXKzUADt5ZJZZJiwei3vuf6e57ZjC4UwTSM1iqQKv49MLFMc4/nnyegzzOX2k3b
7fK03rtfHcNhq0J9rABSDjYBSjbMA5Eltr8KKPoXfY9WFOTSVGPqx7tLOxK/TC3ZSh6faWc+i4hG
YkUQIfcrxpTzclDIpwG2JWjr1PhPWeralPLjc8i4Y136+5nQsfifeK6XhNmbCYpbQJVnzDnObIeH
aou5SCP87a9Z8V5pPo2A0QIWsUtm/D/oGjYwjlOSBY2zQ6b+6T119ouo8OlTtckurxEqNCvBgEb2
q6oWvIwy5Rhli9093v2tszX+DvwiyXJ9D3ft54kqmndHMtdPDX7UWTTfmpHBv5pyrnXpP3pKMK/Z
8lUtMokkzzZqWpHqWEkz2SVyZqwX4k8fSPsSgjeIQtOpBYxAnj1PtXeVxhcK3HQuBM2w2+uKyxKA
NqJCrxZjhgDZEknISdXkNcvJptksktiSMR9bDBgg9OvZ/egDY+//Hd9baE+XKkPaH1+3WHJtTPgp
5uZxfvjAH3HKH3m+lRvrnQSu4yYjyaIBLlTUDZRP21zTIL9g+qU/+vaks1bG8kauwSZL5PFbAigB
2ndaF1iZlz+DmiV+OCLyC02oEYPx36ZByvo2raeFTsBYh01kVlDNhBZld8RbsKWvkmS887zldFCQ
x31ETGSOZgaKsKFu8ME//7u81UgJ7xNygCP2lJYlrif6A5RTK3YjGbBMMC3yQlyBnZRAO7hfVJ0Q
V+dCs9uUwLabU2mCC6XL2lfFEsQS64Nfizknn091xxVeDAM2Jo4wLaw9clq41FJDH4W8DxGjP6pG
S72CxSLQ81inB7tn8II4Yo4Wv1/itA2D02vOuPwzHoU3QTzqTwftbEenk1QKavJclpEe2V3xi38X
X2l3FFvk6huFufOCawPR6GzljXyjJQvHN9gaj3+MNsGkb5A9y0Mj09Yuw7zR7a16gNzGUFNDWFXV
yGh4IXtbO0PoFMaYUrYEsj4vti4gMmTBqHB7P1+qjEKNvDIhQm/sYGG9iYVZMREx2pLRn1GQDiqP
MzknwrYww8sc1DzyiJwdnZXkcaZZiPvGklZOHAaSMyeXgEbA7JOvdfEcR6WZsT0rRozkH0dpAWGu
sAhhkDDN6fKo28GQQ86vyz7kgPXSIS+3++s5e8YCIZ3IZaQLFQnmkVDdkWwiSPwvmeGwOCEbm5dY
t3ezIsYYUqscqd8Brrxa3DtA+AO4SmdFy+P6wRWk5g99fehj8m6GGhDE0P16dOcAU0faiofAtnn7
I6O1S42+wSMdgJGOiE/wL2SFNV8o1oWb3kMrsIa627wRlEfBGL0isShxiZBCtfAtWxWgtIrnQMbR
XVpGDrFrAJDg2SJycWto7uGf6mKsTX3wlYmKM/BlXLqXBDxkSo8M14K70zEfzYlhBeTBuMX8e3yf
z8l3NJ/Rhv9QRObeN4GjdBIYeHyimUkDz1ZUuIsMhmy5csXQWEjPa4NyORDyS+18r1HUszN9dOFH
9Tyx78lSKyKN2niYiy29lHaGu08wdVUjqcg1v4dhn6LL8br+slJH3EtzXCaapgWSLXmksLHYjuVp
z515IwdILzw3XpxhAIpwbxkA0CKOXg2XVDm4B+v3DvIMzQXGxPlqv4DXxeRKRc3DOSf3LsSrW9jS
QtdXXuifzxP2QMHVFYTxNZUnM03D4fQxf63q5PbagOWKDY01J+Zd/uJp9Ktlq1SVZ6tRMEQIqCHu
9xNz47i70gjtpoT3Do2Gptw450PUNEqLz4xdUiuwPEa/6vIb0Xb+a6aG90xdZlvyi46xRKhtX8G+
oAs6rUOcZF/OYWoE2O1fZWkQFk12CPt2zkV1VjbuT0ruUB2D9UPe/NnJCYmBl/jDV2dEsv60JRpE
S48wpMULKusLftrOyxYpomnO3H+DY8lxhlEPVYz27qLU0cDFjlXGqHkxapawCh2cFDWW2cu1GKIG
EaVE6cMMklkYHBbGbPeuFHR6gNoYKuGm8Qm5KvTXxnau/j9+Ua7Xh+Y7GmT+nraiv+RYQXVwyLFt
SqD4UufYsruvr3FgWsTisFxNjUO9UCt2ZbZFBJrIzrFATlMnC8U847PUUDQYCz5q2QkCvcw/zD5V
pNQWA2yJvTDyGPQJgmVHdgmac+YQ64roLm3ZOqZgZ9Ha8DBhlvpQf3pqKEcGRJAU3NQOsxDTrnEf
j30M4KEZd2bXTrILZ7ITbf4PX42qZ71aGZpXIt+PDJUWCTsYIBYxH3Lg0LnNCsPARU4in1je2u0g
j/Ttcmtz9sBPwa9heQXHN3vBzZSIIExPlTLCcCevo2iruKm8ojy3OsSBN4vRYatVlEVXND002dGf
Nqglq0JnqiKtaFDwzDMzjlmCXLpnVDIK4TxPUFa+duKdgzTEGQICqiG/10WwjTtqgXskkdt1ANcJ
plAgJE8qpochvDW+2HlWbgpsxrJjeo4tQdMizSQF0LbBMqgtbG1oXue7t5iNZfQCpuC97XN1/WYo
J7V/2ShWkoyh28bSh9jf6naNwss4Gj5hqXpZD2jyFZK0C9G1WBrCMNp2TEDkkDp6u8qNoQJCvEtv
kO/tldYEl2hTv6mpncQey9pMf+OTjkMxZ/6JFoUeyA12wxYg4tYNTclnhme/qrpV6TNHbTbYb0tx
ba3L16/RTTVGheVuHq1dzqmp5PdN7QPrYPUbfD1ISSUuzUVK7pwjjuSRViNi+3l5L1BxUBMgvITh
5G1EUInxS8RzxKsXTHmlk1U6qKAoOLV0GEZ8CAMFK1mDzjKoClLaMFq/8ZL5nxT7m4d7URMN9tXf
3HCVEau2B2gyU3gfTN17NrCLuOAysNBSJ4xCgz6P0+bQcmcEbJJovMGtlGZ8rhnmY4HecaPR2F09
a0pW8aV36YBEgAgblFbQ4zRIVVezZTlzMhtWavfEooHHfquVU+XpPtSouX7uJImBVd0vJZZCKtDo
0T/QKyLC+CGKbwXus85Nbn71R9/+TJ5UstJmk7szV8xgx77a7289gTj0LTohli3BugAJ56vHm/e+
od82dCGmMk/KzkrJoxhxI3XZYbZf3GWcr25OcJ0TMGHoa589RokQm1KzaxcvMHhDXQRwE4/JaPhc
8qUHDDNWl/u9ZcDOXEd7UQXnw+so0E68RSKR/4RarFb373ffNkoN6YIrRM7z0qufHwfe70iv0ZBJ
9+gTFbW0UdvyH2jPQg3wvl6XvFIKm6Op+s2K3b+ZVf9ImZKYaZAZTmudmn9Vj3cexmxmjrt8mnUG
Hk/KoqH7RO7fU4q5HawbLu0iccsm9j6czm5dfPHRfCakY/7H11ohocoOHvfW/DHplFLMf8hB5mQi
7KW1A10rIi8xVv1z7I9KLPBPKciaW2QyT/xVfO+VGYBwZoMr4C+alN4UxUcmbHLgpwlwASKSflp/
MQuClTJlc7X5K+4+KsqAEQN/dkNxvgupDY01nNZnWdeXTzhgWq/J86VcDkJVRNMda5uaKbziD9ay
Z+ZcbaUSLDozBMBCnshjTWwodTalYpkixyDAkgOpCBjy0/ZebrKUK0yjWpY4mzqKBttrLnbr1fXv
2B31ULayN5tQKge5QtnJ0nP5GDCJcgckgZyDFT8/98E2vM3DmOXYn9COI5+WbhIny+E6LBWbVikZ
6fbyxwvFrto8mKrMpo6SWfey5nF2Y19O2rOpC/GtIqNvugx+0qRttHZDxM+zHlOS+s3prIb3FOgX
MCL41XE02NT7NMWCbEbXlWl8qSwNGvg4KWTEP0/lUGmZo8Bbz5hYehezh+iRqPJfMmmos8AJpEfC
CJLnVLzd5sNjnPDLZA819it69cUw+JNrt/4t053xSYmdp+zOZ0RBVW/SBobMHuI8Gw7FJZd1/ZJJ
rrXtTgiUiba5/4GU5tf3sX66WTaHvC3TCxdYhDqwjYLA8QmdWcl6jAiYg9TViCrHOO0/+f2ePN47
2seGpZpz3iu9ZfJz5NnZKfRQBJnP36xpewVS9Oret3SOOcctoy1BrXJ/jrOHTgtw6/J5gZEpUQrY
RKg3A2V9LQoTsc+bXrm+9M4BfU+0VeA+ppKMCaRSwG6Bi39WaC08Bn34sfOnS+AL2c1xRc1WKz+O
rMHBLuUtYO4oyCINOzqpBVgFZQ52SIhIpBJNZaW1y4sDIDjuUeoxlKZjfALoBbJ/FV/EzbaejUrc
Hkq9R1WU+jZwYm9kAt6+1qPXARy3mj7teDcxHyZjLr8oKIPkXXM8t1FDnU8EJpM0gtNb+ceoc7M5
zQn+gLMEjh+duNt6jDb1gHGmu/KVmMkmxUbay5w0bsnwF9G9J/cenL1B/GsiUeetjly0uyFhvO72
8y+DgcKhShWnZ8h6OgGczv7zONI4gK7cGQjJjXLQSWZLFXNVqIZOYVBABgjBeC2h2MZA29elcOi8
fs1kiD5MzSAaMFRYl7HHpdLNaqYDCiPD67nk/SHaa0BWbzeLxIi41oQnWN7kIT/1kbEZGQJWKLeE
uUD/19VnESLtVLcF5Mjnm0Y2TuYFWM2L+1iZmUidwgVZTt925btPu2KlLUHC1rsQodqiHpvkuHbM
lLhiXikL2dLIT8WL+EF9BRzoD0UQ5gBm+pfnhN01V/wUpGQfhpwGdqFPVdp11joa7AFaXZRXCxUZ
1GsqSrbXRwRp6ndr+59QM2/Q+0DuFYSVZaOSt/zvME6BbnR3JQubzk1QIc+35puUKn+sxqUvfN2i
VZ/MoVkkGT3oY5Aw5nM//NggXpCkVV1GCzh1cSWjRlwi7aJG7vkr2+M+rMf9Em8w47m56iaOgDLI
j2TBCE0EC438Qycf0mK/msRJVqE7K8uiUv3cCJd/lHIpbxe5XBFsk+DNmKRR7wTHfd/JxFm9lN1L
KoLtBZVst06VUbTc6AMOHXcymD0JqYdjvm7T+UXMzGdwz1oPYS0QV5WSixFxlM9PU2fAzbqPFtcr
IlEJLFFpZHWpLW9yvoUykb2gGurhRtHcxzbaZ3w6urhTKfcy0q+U5HJAF4103u92ZkVDtEyGagaS
UST6Ya8Ys4S1pDubjszoWkJxfUxD8LLfS19+XohrXkzXQbr6tXrgm+sMdevOtEjfGysv3Ho7EAdq
JXLpl0CcpG7TYZ8+FuHnMkNFlOZ/kbCgZ5UJ/B4VXaKW7eivHNOkt85GlpDLmsQ06uiNPfmGgdIS
3C7MfdB+zNPG/57WsGWbRkoon9d54PrExicgczHhpcR+V+hYqFf8eHgVHgXnvzEM6bw/gbh6uX4h
enBaG/mG6CtCIn26DfMXCaE9Bz3BtA1toGTFEiK/hDefkx8yAH4KO79san3CL1R9ImpOguWWqjoY
JQTPhxleW+l1/0TpS3ZKGnboLt0GvSiclNSmORjBtXm3OhNKxirZjNfRegs9zWz/3genwbyTlnOA
tUv+7OmckAq1e/l7i/eZ5UdkFNaZrFdvK3RYaLdbBySE2SM8/QVbt716D+jR0G912nmPc6tuntP6
m7Hqulow3t3ctYFcupKkrWNiyoMWuNp3GnVgAuvgtjvoETQiEi9085d/5WtWaLc99eZg6qOVjlNv
kMP5F3G9VpMU58/wTbx3VKmHMRDzLwoOwMIrsWBdgT4QAFgEZbR86/pEGZndPSWvvzUDf7ePi+Z/
cyHWD8zrdrus05/AlPh4IkqGRKz8YLooi27dnsIEvewMazXp+POONaXJ/hLFDK+m0AmLOJwF16UC
zcbCHZCFqEroG+br7ASGN/o9NYkl0ccctQqbas8eIk56f6ij7qb22jcu/cNTU68UXe/O4v3Hj76A
oBiuTEinK1051vXK5QbOySvuUrUd2OKHETjNIkm2r7jeuMKtpWu3skDNbjnhwbv7DPI+kYdZAtZJ
j/+pYK5eb0T5P+4gfq8l4Bx9FM4j8z6nN45z74v+dRtAnodGVnra9Pe7vWQfLoIyhi8iPMUJAE+e
GJBfmqyOknqqamqaP7GaBP40Z7g1RdporG6DlNjkigj+ZvuTAnXpVPRASn78OoL5lsuJ7tuFsZV7
C/FV/zwWv9vExmTt/gmmqi3RUCYUBphySVmHagh58wC95t+By0RjOx70W9xUdxqIfeim9CDoHARS
XfXjlrMVOHFGpiSY7pKR0S9TU0yHRR7djC96bDWjuuLe6TKO9u39ITV++v9uSvkMJfw+HsJG45EY
g19LuqlsIDUmDiPHkOwQYerTWS6whDtScUOyZ6OVhaYw6BAUwYmFyHX//J56MHg2K/aOfcyjh/Ck
bF+DnbpQ4nZmKi1N0eMdlX553gyY+938WDAXau5B4u09ocQMj6E8taKCLBi5Y1p3b90UGO3cdp3k
iWiDWiI3hUCddw3Sgh3fdMNYWSlKiSiK9nM2WBvIIQ5GLPK25E2YcyipPnx0Sy7YGYRvhUWLGNCu
seX8hX+130s75hIXq8mnLUhOREzr2UtorT2uzETHJowepmcfPdaSgHy5RHxnG7qO2AO67cwNXiHb
C6Ly4cl4gx/06wEExoUW5F0z8K4LQtvdJAkYW0hhX5+VcXmpi1vC0PYOAQewL2ctkWjueLqJ+ShE
CQ1wIIUZ0nAkjq4uqNNW+5fgg7NjRMk5SH/gANGaIER3el5/xX6s4EaNeuZnNPwa1wK4Sfjcm7dK
g4u7WK0jizykcPEdJ+D2rcl6B7IX4MFcPaQsf3yV4F4LTbv0LYReI+M51F8z8iKF4+vN7YN0FwPv
uMn0KRIQ5aIH77tUpy6kOkk4foAPwDBfqxUay3Tk+gEQVgB0uIyZSzDOmibDEI9qj6LGtYuG8Qd3
xAIBP5m3y5jLai0q61YPb04ENNY8g2U45K9t7zyWabjpY2WXfEzgnBYV+qta7GzQO61ElP4s1yyj
SLkD6OHLpfxGwkrWiiq2aq497bHY+GAp+uwRvgSUiYE5Ko2ewK8efMp7TGYf9IFt2xSPfsRQhOZE
EBrFIHfND9BpUNCgFUaQW+G8oV4f3kT1eQYPHtdtkb/1fLf2hxAFa62FKG8cZoUThY2jHILkR291
WqUcTOrPeoE7uPtU1KWuG7yZiMw2zVoXp4UjVG5oStaT4UkVO4WtDlUbNgXZZnguK1Z/+Ty8O0cj
MQPAVL+YmO3zfOX8i9Sbiu1LUzwshOzvOrRiN27tvFD4BXjnzXsVwqsLErXqDQ79TfbFOgG3Fc0e
g9R9eiEGdwkx6HVXoopesryG6d/pRaY0l3s8nRnyWFGiync1wi0Pydok5uru1jJUPwSGSIUhPxUH
msE9bofE8lIeraL3pMnErv9RLwFA5loF4Y0WM8wlSJi16Kcmf5MnZiuYNLRm0lxLZnh5rSKewqP7
Si+hUH0vXPXaAnQpty2Qr6+vr/LDxnr3U3x3hhxhA1Q7HJb2okjyfLsptR3ANNgZc8aHY93DWhcL
qCTK1QU9xQDgNf77JisKGlEqf7mhbmmPyQygnuDyBlTNFRph4Gc0Hao57Neg/hqPo9yJag4SP2sV
k990FCCUx02xLtM8Nj3JehyOr6tcXgZSGe0sqQDQRq9/jZhcqtD5JH8RM7R4Fbouscq2IbLc81Nq
b7etvpjpU04tugHDdAgqD3sass/He/+tCz8ZRtDb91g65Kv0KTZPYy8iij1nVmtrQBwoRG2J88wF
nEroS14ogKTJNjKTUrya8Y4hLITKC3AuUttC2IwLQEjY7je8OpAwzAEWaatTd1DKSKraYl55HHTh
Crf+JbXZhe8jhx2guQGv0QvxgQeQKvCbpgSarkCadE78b0QIU01/hI+ZjsNEv71ZTPgknDdJmn1E
c4BJbxwMlKpsx4UtvDXcjXhJeOD6yX7AUaRgFt7hA08Kvq8devJVh011Cj7GD6wvbUVJlK5oafdM
SzCmCNJrRpYdAt7N+OEah2u0qyeKeqSRQakTMOrwxhQweCe0X07AWKBOhVLQ1p6AkCNyLEh7GO7p
NJxin57cDH462Q3fCMD5RUOtuti1BR/sIZcjQKHa6AFZJYgU1Fhu+jm1TZsiazRkCpuIKYu/02NR
wvCT0kajPGhn5wI6N6TfSED0Ox00hGVzygAPSKYNcyVWv2vqRNnHTPPGfX1xLZoQuoa/4+Nw30zw
Ch3Zgz0Q86i5xsHsiZQaLGyd/0Ntw1BShxxBG7g2VIosT3wX0VAJlCuBGhDPCKsZBGoD4mwRiEeo
37CvI2fp8+3mp0phA3qTqDONxJ79gPALGTvSR/M0ADLozRku2eboqhgIrrwG6lCYeEmb3mEsC32W
ZjI/DN3ZXrufLEBcaDKTyQYmhaSfDtkj02VZot4/HFVg6I3a4KPMCERwL1MdzyPqR7/npdOCZ3oV
k104txftbi5KkiW9rZndrvGitm9sbLyRaB08eoQJ0P0sCSQd8/fHwMWNQZpYDQ444gBC0jCe6bmB
FwLY1Li+2Qy/+6mJMf7SsIz6p4aSJlBK49RO14V4xhm9XAPkrfuV5iCTHtReKzgzKHMFwtL/5ycj
w26WNWRQ9O51wIV3jbhrYcV2+Vjy0EvvJBkcq5TejWtQK37HHendXcHPlvFJSIqVfSk8ZN1Q+v9Y
jnp8o+AiWsyuVr7oYJYaonIEmh3tl9q9+Cz1Str6qaO2cD9G7/0hCmn24aGup5tUV8z4oPX0gj64
z0zICDSGbpHNsrx4W8yTNPK57lvEmPWODBWNwmlOWeyL57/8ctJS3ANDW9NM2+Jjap54mveouN+f
lT9Mr+8/DZScyNRT95JyBw8hAWWHIFJzqp03SO/XTmIcc52WRVx9hq1pLBT2RUt9sS6NZlz0gKH5
VKTNNeSog/EcyFnxrU8JUKeYTIznyf7QxIEhEa+dqudjqzAVyjjMFCk098MjsJ8BUzJA+nWhIlEJ
D8rAXzP1TZFKzb9up+at4Q1YjbhfHNkt/f8yDX/2AY8h2c1ErdFr0d94bVFUyB+VFUKG9oBQQk4T
dOdfdc6wzAlImBA4oBX9nkMZYCHDO6+Z/Tzs8W1TbC8VEynuTEfDfo3YM825rdylqUeeLLslnjD5
QVaghe3Vv7wsd0sXtSzE33r9h3ej48IZcN63qaSF6UB4dNXL3XdshJhgVL/WvseyFafDJv47ldkw
NF0H95++7sLf//hq3EVDiwFn7QTR/q5XgvcOuYMlIQ7n8AMZwNhFy58y5J1NDUUhft+N+prbyaML
nn0I1Aqn8B9TVlEsiBHeHfy3bwc9oB4QUzkPXsh48cBBDOdwrqaaxQlHtpexzL7RpPCY7DPDZp5m
W6ShNocnRKb5Dg5b4U43jNDFSwAC4ovA97v280ao8Aj6sc5pmzcmXyQhJwbCXqS0BleN63JTwoeW
SOHLU05VmXX5AsRDPTHLLEVyba4tOMhDpbJpUBco0/20vLN5OG4r7YhuBQsxYg4ulbha+KErF4jE
mc9+rBnOvLPH4ecfFTU+8d9F0XeqIakCZdmb92YHuTMvGi/sO6tFQ4aDTtZY2radgUHot7UPVY53
Z8BZvq+biaQUNFEbWrdUx4t0+dJ/E4ozeOw+K8DMQkcauvEnuDhkGuXV9200/U2JPvzb0U1HgIpP
SnGR6c1+TxnfKxyqbOZdx0gjnMMhgtKuN050sWxdhAdugvx1KSNbB3hhsiGP10eSDNhH/ymefEt7
+FFcSupJzCsO6+HU82B/tkpv8FQKQLrfMlVE944uecsSg5sBQZZJdG6UPQiVYWLqzRo+apESAizI
NlnqlKw9HV5rRSOHEkDr4Z7PZDXG+EDfOucxcoWGPz2CWGi9r72Q5ufJxiV4/NoCPviS7CGmYXOV
fwFp6J1DRcvBPz7SAzU2hce/ib2iSt0Y7r3geq3+shh+l3eWCMFs6tRK3L1tcR5iWQkLZeCa7fsx
n8lkE+RMms+Z5hjzZBOPIMW4qfh3i+E44+19Linci6bMacSIItVBeRzVH39t6NyfjxhrQA4ge/fB
vHK0AagewCT03ezqzxm0mDh0m40/CeaMcWnDVJSzGYJYEPQ5d9Bfh9APQ34HnyQrGMdwoDbus2s2
nseMTK9y+gYKvlCF6SKF5bCZa68MjMllkBniULCxM80IB+WCyFwIOiMVmwgruR+fd9lUZZSLV3zT
x53LgpBbuT65ju/8A/1kDBvO4CAeLMppFAxvDd9dqmqXVe4508LwW97wgDyC/L0yEGfSTLcyJGvj
t+lfSst8ZgLRFjsr+KhEahWbpZZdsE0Dq3sLQNgtuavMfoWZi5bMUu1Rs/vGragz/Ykl3LJrpOla
oIRZfwuOSeSpKY9LDH9uY1dwCYNfn++vNQn744rxyh8u6q3bVaZ0RZYc2R1d8T10M8c4om2mJ+8y
E5TYhJm1G55hBgl5pWZgs/k3qiGiDlWAVBhCWZ6TxnKHtCytit5T+gXf1irxxnT6skRRSaa+T5rC
IMLj4Tna9eZq3FSl0VCdwg0G9FRrp6KFPCf1usV1PMxeQhP4n0dgeSiBVqJe9azrwBsQHw5xpe3e
ReENsl/X+8yLf6AbgDvsmA6GwwEbw/aSZkUuXnvLL56nVJBmXj3E/H8ve38IfkkNTBE2dew2YTjW
XUCILgnQj9lhcCDbt1u78INuEDDy0U3rJLzaVtfvFZ7ANGlZEzY0ymO7ZcVFv6JKVfdGBMHHTXn1
nfGRuEY+Pg7n3629I7fKJAwsK5Rq8rwQue5+SVlajrw8UXJpMct9+/itCR5/eoD1G+homGRh1nFM
4BDApqQs+0hnBK+i77jSVSh3ZjLparIC8l5X9t0N2VJRGrapFZVBVv7orpVbm7rU+cGOdUmwfpm2
uK7KKz2v9a+chWLoz5hD9QenXVkhB/NBX1RvJ58k6ujb1+SNhsoTGaMbpF7Cv8owrZlTxzcuo908
5iGZkr/E4GfGjBrWl9o1NRcYn3KqjxVf9HntyWRU5T6D54HyE/zaNaPhBW9dY89AwxwRyQkeMhjV
/vPNZMJY+d0Gl8Em+pU8EUUPx/Qj1a5tsuzcEy9LE0f7y1JOzqY/kuiitf5wUcH/OyGTk35T6ldZ
pO5vOmpox5H7OMoDcSyIscl0zpx7eokr681J1gyTyZ6rMV6/p2FeNm8PxczVH2vXQOCCaIeDuWOM
x2Yesqz0q2VWuj+PRbr00GDFsRUClVCkIVKsMvpiM7JTUc1jVnAj6iOktbqZeIJWthexHOEtKU0F
ZOA4WUrlZgasfuuRqL4ims2k+Y9r0LAZc44jaMHKA1uS89127q9gnDaa9tUmvr36ndM885g3pJ/r
CyNVng6bFh81dHXSsr0vI4AwUg2nJUALby1vp/fHQKiD9NZKS7q1mdQ5aPk4ADHrl1mSAIJrmIAB
uQwLZV8ViJvnTu+ljO66gqW1eBJ2nGxW/dcjQsQSEzTYsAbAuTvV0MCMM5i+vyI5UJzeITTDY/CN
Ke23Dh9qHHUYah7KdjIeRvsf0xRnldbXOTClhbOwlSiWyj38eO+bsiPwUxGflP8KEUzZi+9jfxRW
+C3rJ1UpfXzkLv4H0Ui4TF3Fc6iLCsq8+b3ZvXMAAN74tx9o/fIl8Wp7xwbUlV9BvhstJ+ks6suj
gQBOdSvXmVY9kOmwT+XJsB6RGpR+lN5WTE1oJGzwog5PgnvN4W1rDd/F3eBYz7KVLvJhe3W+V/DJ
euGiWwYPD8Nk/8tzZBTyVndZxRfDPN0Nz9lpqUPZ8XR2b21NWZm2FkOfDDv/BeTWcmhpkRQOz/34
6estd97yeOWkQdVh77UQ4s7A9uMMZ5BioedPB9TBnIF7f8dTeIa4+wL9ksMA4DvmW0InTSYEw0Cf
rfPmDftvsGNRRnICwO+Q4+RzkoH6v+vEnVS7sGOwyvNukM1hmP+gRGszcdwnA8rG2HqmGWvWFqLL
6ynJMc6c0LKCnvBp0Zxx15vCFlp8l3reIXlccWxUA8XuXjvwcGtHdWKDJt/D7xuuB6fi5NoZ+xEj
BuxUb3WSQxgeGTGEIHJXWpMHUGaCqhSL4lgwPqudUgUBcnkBa2uqCIID/p+vqBV9Vmci++YgHK/P
Rl4KT5O9ezwV45u5BcOzijy1iBaTc0fmj4/1XmekP5MjEyagqpQg+9KHla4adn3hMqZBtvUXrfIg
c4IeySqaPbHCS87ZO+U/fVV7sSMVh4y7UbcTGb5V6YeVM8Inac92hbhFhl/ynMirWKF226rX2Ye9
pQWoKvB3OOdlBAYy6vmG6sL2r1PC48urXSoOmaNtHR3jJWnbEL9IXQZKLUGJj2VIsztGk09dQsKV
CnY75GMTvuN/Pq2gxmJLysOYU5OLvCI3KqaYMAjpuXN5yF3Bvs2M3Hsseup8DPYeCTpmoAEvrVdT
wsnp6QSTPKu/oMyijns5nExecoo4eL9XaNcUWC/ztvX1oJmbbnYRGnSornbdAkGWz/8lg42EBgp2
F1URttO5BlSdcke53F34ETBrDetmUfJrVEwlhknDBZTFVAh3LSispnN8VJRWRvEh4nrO8UA3swgr
dcwkYQMk3dMRx/0HzK3gcv+d7kPRY43HSISs6JlY6aTGENqhoigsawIer7X7LBUmYOpZhFa5ZrWu
ZmGBDmpjiXqWIw845Jo9JCGHbwT4mSWYxtWnrpWUMr1hSeqnsRQVYLQRqFJhJ4uatTJtyJs7AwZR
gr7FfhMYx5UhRbDcEaJmdkqblgfea2a5GnsLNNDzINLMnHAddu/09FhdfQ289qAC+yVBw8WstlBH
z/sBF02GZ980DbRxI/ocmJoQqcoptxXwoIAO2mfa1LdTIahFna54NRK+iTwXNbKquLQNLl7bfwPu
HKM3F+4ovv9m0wKea34xRd35VYu2cqWpxkLNbKaXPzD9fzlqD5h36XbBGRlrgMai/76Ru38V0pbp
1pDRe42S6u08oJYTjMB6hH3EWswRiCht+rMCDph2TzOFBWGGkmuRIVAyNHKkR5YcNfCrgiRwsjty
npM/dTjxSFrAMHFGT86ncpySgbCVssOkp+VMPEGXwpasezJdY8junMNBRW1dWftBwye3Mwu0MOgT
vXfGqCZ7+7TcvSeH16ikCzNce7FXc80jl1U1bv4bLMoGwxTOPQAy9g57BlyPwtew064AgDdlQY52
Hco6MXH1OsyStjaHM4omXH3jpH4tRdPa7bN01TnXdcLCK7J5VapfdK2ZGi2mxExYuWtSEuxtNprE
p9u7hTjnvN6hCbSAmzXA6/AlmUNm6UHuKoQNTPhLPFRvgIMu7oKgiZB55bUt6zSn1UdIh9eia+tL
emFJ1VJXx87Eq+AnqYn8riS0LsGo7/pdL/lYvj/CDl3U7ZVf1KmTf1jg9smrzzkOOr+FzvwJkAuC
f3Q6t7G1FANjvDpwE8O1s6FiuYRYCQHSGULBB/XxusTnBHrS5aCOgmLNgZ1YIE/dupJ2A2PsKn9m
xM+Fmq4ovcevxGdfi7b1V8L6+LDU5D3qghSOr86/SCzd5gv2VTnn1MkPyse6cMevc0pnqpF2Ytdl
sYcpCyHfe5RcbQ9Mk2X5byLdhUMVYBunbu3HyDkppmihSPSnb7LhOugBVK86dorYs8z07F8mCH3m
Lbu0I8NRl6vTAI+rZstt6SsW8XBBKy7KO76ybkLH83K6gyd42RWJmZCC5h8rVFYBDvdMws05GGM2
7okNYyeehOhhbBdbb3K2lCyF8MQNn1bfkvjfJlckZI7/KXn69C/RMuB7RaFdT66mG1vfyUPKqzzj
scJACYocLkqsiiBOcjD74qgO6SBC1BdW/D0gIfST9zQQAO5+8/qPnEWhPBGU3Hf/2cWPZ90VDjJ0
UBpDDvXByZDClS0xnjvAK/Q/tXaXWyvE5oFcmAg3cuJTJcky3/DgENZme0bJCMqnijEwCZD/y3UY
cbx57RQPVr8Upf0/met2xJ8vGdumOZm03OB6/SmdK6uy6IByEdcRGuRRxfaOgV1//LtfpgzhnWlB
GRIxNgYuMHnuQCNgeqrlEVjBWWWzy7jVwj1alPkvp9H9yRgdwNqbL5OIjk9AJUNgAmITuXA1QSEk
hkew3NdPpzadvYV8CSE1dVQp0niQTKZfe2MjaH/jwvU5gaQIj30nkmBZSw6R4YoL4FO2FFQjy13g
W5EUoHeYx+QBbm+SqZsyy3GTI71osUnb2lI7Ue7rz+w2piBb0KSr1sCwAopasNYNMRrZ5qM/p15X
QO2B83ibPxRD0b+p5+/SrIhorY53mRLI3Q9dRoegCwYys0eitLYNMRENdUjrUWMTffY0J83wYGXQ
fEq+mD1uAGIHMLQ3bxcGS2codzqA/gJ8KgQJYauQWmreMyeIQ92JEaiLhCdeWTg8pkeimocrME9E
nH7ztzCl01VIsyPE6iXCxT2ANfQZjvVV9cPqAj7E5Jlna8o4lBQVizMsCAQJtrvw0HEZaO1OXixI
S1cE+JLPFhH1pO59RIw4asOwTZkF5gkvwZ1aWh9NUGc/64uSiGWasCfYif62h7C/w4sfQ4x13yHU
CQvBkLgwr5+omwzOYMjivKBx+UoefsxW+PBBk8eVFEZQEa5PVOnrMWynrlDepaOrL02n9ZcIc5aO
J/cY2kobZiWBkB6jSv4yn5IN6nBAeS3fZdgrm12XXk42Wr9FOm+PClG9sD5Qoji1aoXRZQ3r6WT5
CKNIalDwUeXVzI0D46TsH6RJtdf4SrpJAUChJUVOWtLHlZnZmVSqA0nHdghZNvQYCmeWFk6U7IhL
a0DEdyE+V7xx2dfLD6gdLTLo2q/1NaqS/RSZWPRIAq3KMFadVP0rpmmNdOzVZsKV/OAsrDuGiXBJ
bLgcyEKokDyzI5x2ukvkzmJv52ljz8Q76taPBMVtOw6T8shMNONP9JzqbC2Yh5F8gDY+nSEezYlU
8wxQyOCbuoJmL9DhsZkhNzD8FlkoqkPjQkOMjQZ0Zz54eSSPOswmjMkaK3BJI/Ru07Mrnbu6OwaR
LqJmD4iRRvqHkpdx94YW2BvQFqpfupiU76dzYJ9Y6ituoOZQmpl945CntuMGEtsSlYBY433zhQSP
fG6+t3RxOrlZ9ZPaoKlu4dnUHgpcG7ECKjsl4cFS8iWRMRRCOVIYF8Psjckp6X6NaRPlgy5sLjHT
X/7jfzjp2VqgjwsomIg6WCdRcnP/rfWMYXusDXdZBNS35E/4s+Jhm1gMVN/NnLItG6ARtsIQIDdn
QpYWi/93hlrxNwnAGRV8fvCJOKENY5QBdX62o9wc/Nn3rJ0HjA53LsGE1YwEebOu9qpPKUDbR5Rq
PnXy0usUBbX+4EcHvxknmpF8s7M5yXZDQbsjBV2dtfQuEeZWJIKu4iOMuafrMjnaU0LQpz++GRVG
PQqWMvylEJkWd3ouukn62cvXDquh9fdOzAiIsRta6aXnAgDj/qy3KemHGBwAbHJ6vIl9ARx/F79/
nBrc5jOxiJr+CW3DDZ4hE1v21wILLS94ZO7eTylgjwwEGN1kR+2O6HJBAEPXsyAWWUyBvDrf6bOG
r5l1uKcdMnXw/JLdBA1pRnEL5QJLslIfvy0oF+actP9ufu7XmBMFbLeMUzM+uiMV3O/ts4yhYEwT
8BHm7MSLVv1B8LN0oeDIwgwKOESBxn4zvD2bR2kqpM4B2wNkmRna5wsh1MXvoGaTuxqF9xJX8fQc
U3NQcvUZP2qe4IlvFp+5NNBqzRsKcfJ+xtxRGLFg98fU32454zeUujtjg3c8mxv8q76cRH1BwHWD
NLomZelp7pmoAlD/uhGaTHp03USHdTczvPcAp/AmdBPUDoyobcYrbNvwgdIafhTsrvIEp1KxZ76B
IWOOo25nW9HjtaMJZ3dh1C4txL01BW3e3q8JHeYKbsNA6YjA6gVtqW+bSJMLsNAYuXyGz6C7G2VP
w+LZ/5witXFg5AFD9SS7TNpm7M5NMmyd6XBYW+73OMc4mpj/zvXKb/c3XvzLa0sqbTlceOZWYFHW
LcqB8zv1rHNJ5enKyBPnguV98auMIVn2cHFyYhXinm9ynaTIkG9+0oYOiIRseMHp2JOWQgcHiql8
CTWcIsnmenmQLFiuy2Yxv/0fonarxMoZG4OYD7vI5HEv3pBX3Cd7rrgezAp5gng4Y5FtEURfxUzp
BUdqLsBv1nTIMZMbNSNElFo5/u+W1KbETr6YnEsysY4yrUNxJcugqOg98tlg+fGlAOEG1kZrrHHm
zTHK9LN+zaQGUnQv1ZXg0y+2EKyE8mjOQJVSqoIZ/nukBG/mXHattdfKH4IFyB9KyDCAGWKuLEvf
1lC5qxgLViSMrHjpbD2NkePVI43gN0T1aQn0iusKXXk1hK/ZHkNiW09juCf4Zs6BB07iCB5+0gWi
fpQ8pX00sTPjrlPLDQkPf81bxdvXJtAPs/D3zV144E/P0LyBkOvZP9T5NdgVKoHk6gQZgrUsnLyt
3qDd9B3hTBE/3K39FKL9Fgqdr2SEBpg1wok0/0MEyC82RS9QGxMXSLIAU8FOQX9oW8jOUAvtfu+8
WP2uzKRxCf5IaiX9o0lScGtSKSKqKaROuwt75R1mCrqFyt+DCJGjwrjibTh04RHpcWXkizzOfk/W
/nMWVb3AVgTU8mHIDIu2aUyHS1p4DmthhZvWxKJKaIJJM3k/VTsWaFB/t6tNWlOqPjJdI3p1Kv+6
dVqKDF/i0NCEw5KW5HCzf0N61vgS1DMxiVNnf7BdxdWQGaarNu9sRx6CQE5yuBOxm3hIrqQpybHv
1dknplsUAp4NKhBzVa+rOKLRDRCG1HEsr8ZENeUwq4y1jxJR1UPJWC5AqLZFhvJwfHznXhiTTdWh
AJkCZ4jMNymBbiUUCgoQuffwiIZVGAtonlPPAhN3vUDrlkH5phD5YML0W8IUxWARnbDiQughmh2c
ly/4Em7x1xTkCNc+/KSEPpatv5KGt5VKH7LjlqDBhdFXTA0vg4XFWewGVFOkyZvzyspTfFzhwsEb
bsgHYhPxrkbAZcFYFOwPTYuKOWTyFPz+ZHL8PTLPxkaoUNaCNkrgQX2R3OIBQ3dkACEAWcv7Enzc
dCV+oUZ8kaPDFNDD4GisY6nwx4hwcGkFisjbRODdG9tu14yQo9kxU8u/i0ZNWFeZU+PeGotNZd/O
kfT/j++0w/oLEiQiCvShPrVAdFnSevZPWM5lQpuY1k5ZKzHr0sVWgTTeUGLETSdMKHb4wjV+PreM
CzJ4r6s7Sd8HTSsdT2oFPFSY2xYDajJErZT7DY6coT5JMsC+m8UycInNXcUXWZ3+7ttoQP2LvjP3
VCx2ZthzFzsvmcdnwXCqJsPsYbpWPPIU+rmnzer4rnFRVJnsddEWnb/AfmPkR/Z2J6Q/N/7GQHnG
1kBReZqvWPJwscbth5VpeDUYNmF0+bamj7CHhsq05i8wIbK581zoCEB4qDxdBKCawyn4UpoJk5KH
+CmeDEMhW0OEat1mJMKHWCNvznq6fyD3uOO6n5Ji6KO8KulgcBMxBo8cNo2WSxfL+yMuS73cKd9O
7XhRUKbQvmCPvcIV95M5j+poNA/YYK+BcSx46sqTHNEgn1/MEtbNuGBM5K3cWf9FVdZHFCSjbBST
58N5JWBHqyu+eHUuqrcbzVAxDY/eYwk/akKC63A8pZXxtAs5KQT39i8fHnieG20CDyGhVByerAbl
SAg1mLmjGWqv822Xr+6RhxC7GPKr5x8/0ZhQBZzqx6UV3lOel5MUD41wTjDynTDmxTDFRZLp3nxP
KzFM2GXvFVsX/ZVMYV3HkdDiscKXCaQiAKwno1pFSYuDIlUgXQhmCL3dW8os2LYoNzU1yBBctSvt
m5OLhPiOgb8BwrRH1nDptAgGm3fDM6pVVAJofxvkXmj5wGImyGNuK9nT95S6f9xlbLnyyNSW7msn
eWf8JCt0d4rzOHHUDk+WqK8ruY79M1VAoypISZfHbSyb4Ap3v9IiESfkz6XnQfKM4g8kxWBWWBwf
9mFqV03aLolKCgMVtANz+F3l+UFcF3wBTL1cbjAriZy0+8c0VFsmz6u/oy9G0SlELjy6+9b9OSOd
Mgqao0Nge/c8vMbwpqHbQqjPAMmAuPAKNERa2PLF4YqChGg0Ny40xNcJFd/Csgs99DB9DYq+L3oZ
TIXhfvrIdqDlkgDod4togSVp04HVF+YmV63Df2HDNaN06Sq9nb8ZfoBFiaB6VHDaaGAu6yds8fdP
0pZkZMpKd+oMTLEVcce1jm+sl7Hq2YIC9nOz/tkyAYVE+61gA4zhwsTncosDWPt/HHmMEvg7e08x
seWnZxyYh8rIm5sC0K9orGqtXRKmTlEMlPRfPYX0V8yhB0c689v4RTketkMAnloD7QCxLeksxNWW
6KOwbKVJMEUZbMJZpDitq5MBHph2EpyLQ6EXHmDUihbWPQ9/d2OGO6i09+/H/rDEK0/28T4qoaa0
H8nMcYYpTvw3Nc/fmh9ISbWBJihojviYFSLBVunwCM8Eri3sGOmnW83vyHWSck5Ja/KjbyvsctbC
Trw63F/ly8SLAe6+9aRBh1KC/+av6rE+NzAn2zI3TjfIc104tATlgkHzLPAoGnnwcGXYHpE08+6O
ndOOGUoMV5Xlt4TnFqKLzcFmUDo1yjU4if1CGPv8RgpSUDiGnsI6UGO9RO5AGSm198vINbOrnLIv
Uti/C7w69yTPmmZJ3fsSbeAb6OsJDGV0Z06qUjp7qTXmXyJaYzyhwnu93vVOa3JIN1m4qKpxFH7T
iShrBSGn/kV2835ZPzLtWOgXVsks0iDBMLIhWa0UWvAzTvuMGh/iWtel3dKNfM8sETwKyaorUK29
2/AfkYkwlxb/pA+hOZV/tcKiKMwoVxEpeVpQqdAb69IVGn/fONSAA4Jaxs0zLBja0FKgReWZ2Yqa
GorQKb7mZKUGelfVq1qwhgiVvkeJv7LAXe8G9avXri3IWZb/YvXPOZlkyh9HE4EPoK+twNhARYJS
LxpSVcSWI9ghZJm/cik2eOqIdrYGWb2AL/BXZTv2p+s0Ct9Ac8fDyTjmrHBe3d+T1zdzXoRWhdo9
vpoX/5n5UTdM2Smvm3py7rBu+VC3S4GdAKta1ivnI3EKdCLbMJZZCFTE57eZ5meCvBt91o0WfsbE
pM4MuUXknbCRqIu9WaYODe7tIGbE4Wy1fewAtza1mHMAq8/cMtUvPOSe6ePEIgWyXsgevClfqSwG
eeuj/kpNQhcE+Etl+rmXtMnNHMFaQx1BG9lReYB+df9u/jBRwLRccukrrqXvkQgXMxXkW8ms8CSe
fktJUjrVkJeaBApAlE5QHimuNV86mUxCf8J0lZix4UyM024Kr84qqVbC/EbKqO6air7mhf63jFyD
udKt/aL4sClqT609KHQ/fxdM+rbYAq1oTR8oam9aYQZ6L4MAkbUuw681C/rIATt4cd7tW5vBsTDU
YjejABWUdEG4wTED+fHGvqFbimfsJXsYxMfXg3Ih/SlYiOaDPE9reORrGubD4B36x47at1DUZf28
REo2fHNMDqyxM59W+S9lTCV32MRbLbYuyLVndqt0qZEu6BRTe5Tuede7f/m9b8ZNiUPFXsSMk6V9
Mzc4L3ThkKjF5XP0IudIIpoNVR+4o3h8UGJr/I0K/unhTteH4KgWqfTvKEwnbxWj0uxVmedkNBmA
DYJX8SSL0oTURiElabgILqZJMOb+87JA1xT2l3zMfwa+FsIAUw3nu4J1YayWpZ3cfqFuMZvdo/bj
vl54bLsJKE9ueTSbruFI2DyohceIVdUXPrrJUugjbKFOEsoz+9d9s7UvLYKEmcldTth7PJ7lxAlY
ylJrx3j9upvBnyOOJD+qgiVdOF1vWkUvAkNeCJMNEivcttpIeDq6ciAD07HdDoGOuv0PnT/KAhNh
UO2IKFTfxVTHgn2trs/vHxGuwZhHXGvzea46C4NlyWhzGv9gogQEqdGece3bLVHHeZfJagUdu/MU
EObjRf8z02N+Wa7bVnQ7M0ZwWZt7943AYzmNY0ku9D2We6uIiVvJEqe+7EUCT7anKw8uq7uSXcUg
sh/NCoM4r706YR6qhRSfKGylupZ0myi3c//PuwZgHpi7GjlbLGCO5r+/7slY0gdofjUwvlK6qFfS
Qzt7RmSpIal4M47VPa8JVqgCLka47w2THSMPzjfYyXQ3g9aHSeR5ZHjra8pGZ60dpUNjb69eNEQ8
fudP81TuZ+wSHOMIqLQFgpsqN0Pu0mCJDznWzIXuz3RRrsYbkbcVX9XZZfv9o3s8LaPsRQ0yXcrM
GNJkXFs/od8GIEc90K2OwY8Xrhnjf4h6jQpnqbaaJMQA7gZoMmqMdUInnbRxaTQftIIPOJxhY40A
96k3O3m43CsMBr07Byg2YJFAkez4i2edqEb+Y5RdsDOGWfSA4HyboIHR082Z0S6weP6ltWvZVjhW
PxJsl2YFYbSKfhY9q/epp9ExFvle/CeCFB3pWSCs23ITIKEmWQcMENDC6R4GUU6ohsf/WcA3FSsH
VW0SO2cyGuxZ68eAq9jznSWtjy5W5pdwpFYiKp9xm+6kHF6hwruWrbCwm4k2oPKIG7CXtPybp5ud
k3Kt4+/X6TEl/a3Bc0j9pzyanwKtSj1NYNaZDFFfed8b3DL2HDsBLAwzJ/UuM3qV5RR4xFkx79nX
1vLMc4GhZRN54LTjw4d1x4QsCLPri29mVD7gNvKZ5qKiAwwNhJO+hLMyt7DGytgEEiqDJ9BGYO7d
d+ITz4EaU5lqjbup/pocXmfUr9yy4bu780EW8WZmrBeS6tRZ/UH34kv3ba6X+Z2HJ2RCXXWDB3xg
wmJcEwgjngFzh0JHy4CWVlUhz4NuV0fS+htO8CGW9wsQ4UydrPg/cKniTjKEPms3Jw8XFBMY+G76
Zogx7SYYCeCqsaDniSMDAJjmAC6TR4/62+j2rrOoVnX4mgad5RpKf/BrvzKGiY3F40gvwDvfXgmM
9YBt+K/1b+HDY0Hdqy0R9gnrHLhIZcZFZ10dZ3FqU+zDPsrjAsNI3x3oWgBmxzMKh2Xy0+HeV7Hs
GbBn6gpZmOPCLI096RgChYDhY+j/UUuB+h9TZmx5SoROGV+TtPBIXuQ9rQEqJElH0fPuazAN/1Tg
TRmP+BBI5K/oNKB3GRWU8uvah4E2TymDj+AXbxOad2+G1zdW0052mAI2gegLGdQ4BCRcOWodvXgS
bTj8h+Rko44aJyT0sP4KUX0bmiZgGkfeZjbG0GDPa54pWIxCLuZgj4JBu10Yhsyv7mUC1kBQAc7d
7Jtb43h0QmHq1fHlB8W7H6JXwSdXf99iHVv9JNyGURKW74UYr3Bd0c4esqIXYPbTM0dEbLa54n28
RgKlvnI5Jl4e27Za6mw18CSGfcXvMonPEAzp0PRysIc9UQM1dFaJpVDx1sjX58l9DlPS0AKYG4a0
qHIthfciPN7jNZWPemfj4qJpVlrx93jCUuv0dZUWQkvy+y7ifIXFT3Xc9ax11MjmTuoAixzXI4qZ
olLqjnSRnvCHU+Ljr4dPFmX8PlqBSv3qJxyt/yAYzcMCSiAaFKWk8szOAMAdYOIwYMUOKJJW/OoX
AelyroNDEVCZFiqgeTSIbY1tta/L0CZTLsRl0OmPQWVxHYpTlkxtE+2qXwnOqPlCKOLgP6mTFJ1O
JgFDSCyyydO1jW0/ifqcXX1cTrJCgPCLzf4Gr0X2+5iJf71/k4wC1pj7LF1ynk77EKGM8Z/cBJlD
Vl0HCXQ4Gy0gkqx0XVpU0J8SvEUbnbyqj73CGasxmEOK7PDqHIlXmRwwBXyLyTGOWe+rmWbQeYGp
iCpp6ZHH4nwuqvgBjjDbSRarXXTfbppfw5aVexH2wGlXi0HOw90GTAg0XyBdOfprKlPphG/mSTiM
P2vSLrQL9rVSI74cF8SWgnfCmIkVhGQeMiZ83TD0MPooPJ/Hd0Z9zbIShw2pdTwFCCkJqEEwyEip
lBRk5mrxNuU6QwiANKbz41AM/KF3VBnJ5DCxP4oh1cC08Yk22YNS6QwhnJ4ddoSiU9XLOcgTtShO
Dz1LD6G7NhmZGOXNDcxwU4Lc9dpKi83UDOQ58we3tdHv/cLJ3exZBr6Mlh6fBbGmWsEWmbXApZyq
LnvKfHWBpVK/RIRI9H4N57kqjhlyrzOMt+XzFEzc3SGGFFZeSwb/E6rrowEdI0JWLEyStSgnhDFV
78IoWV1t+ndgVaCtMzwyCtTQ2AhXLkVKtB7Yiwm+5cUh/BwBVRU8Ax48scFmloNEX/eCks4AyAQt
ytr0HJg6YFU6NXgI/Fa3lhwHTO3gfRpeuObvd7F2ObhWa/DIsjB27Tx4/Z6UZqsWgxyFsmeIS7/K
+ysFrk5cZrsY6I4HqquakZx7NKNDa3MhnjoU53RPV63Qqqj/4pWkSUWX4/2goyoUQbkky5akMLrR
xxENJopW4JYSoG/YT9C4lWznG5T/D8Enh1sKSvnc9RTPPwLtZbyTGpfPwO+nk85hRZXmcGb0Janw
yS42/1Ckptyg71lARcs+rNmPlOX1e7xXemJNM9dxEC/SKHqZGw1R8ovQB7JPS144Dps9+KVLcc4K
rZZHgxtQtHzmSVYnbmxFSKdGTGjcd3En5bPd7jIH/nmE0de+cY456vvitAoi0WGVuwU5hDcC6hxg
WLSUX7srHVE5E3N6lhRoAyWmhNXhch6XQKx1U1rQWIYVVlLYDorz54KNGiznVCgZsyz9E4EBYzHT
lbQeouYBtcVXp2C2Fi1MQcDXa7cSqhLaoW0zecksQ2hROS5uKuttk3rooSnvpDfcKEKVAJOob/Fx
Jdb+kqQszi7zOtmI5IbJBtvnc3NpGnHU28uooXfTleFPAOkgqZQx44uPfrElqnScvT5LlkzjvTZU
BA1a2YM9YoJCxsMHHay4pPd5u1xbsEDGQ4J/BpFDxZW6BmFe2wWKjb4Q20iFazadUjppemUJBeFo
q5rb7cTfwlKKejUXaklLoII9rOpwuuJm5n/16PP1GmLhM++ZHctr7WEcDkHT0yiExSUYIfZ/+Aun
Sk2w3dt5751K2RykNv4+sF54CxW2I+3zCIgREuyF17SrI3+76EpOPcDu8JlVLlXvSE1jX3PSUABc
f+sheIJUjBkKZ386tj1EUeAzw1VM4bAFrGl8dOjmmp8DK38IEGoGvXDeXFdbn/2jaPS+x8bCmlQ3
FSZuAoegEGzOVHEbb4afQB/sqQ9dgsFkhE7cf/VVTw9pOZedbx7FSClSnYx/GZqFFfPcU59BqzGU
ZM6ZZW8hsYtsVtXzzJ1Ib0zgst5bK1e/JkuM8imRAGEmUOQjZRLLqzXR/qylhzMH71tiSzmWkKee
UJGigH2NYt4iVZmIzfl5LTTothZfXHU0B0NUhn+0slSkZd5epH7FI+CuUf7OJCYR2Yj5ZgpBS2XV
/DDulOHZtRYjgjsSnmJoNGmPrtLrumI77vqh2xitNI/GhhQPNwST+v3hw/U4dqW/6YGwW0rNNWyB
vvrfdDDcSrNPXiQYzBaFR24on5VOrkcQO5zF5q0QbBp5/eI8Fle8S4Zpap+YfEXZVBUnp+6u4ba6
AzXAStp20X+16ZuWIWDwNPVzEvWflzn9uR+fUKcJykyr8sz+5yfjRazON8KfODwdb7qv0F9+Wr4t
N9uZnsYXJKFQs24tM8vhDBPO1GtnJrnyZ5MzNnnPwhaCyCucxQyNUaCeenrCylPlhxi3pvf1yaRl
c1i9K9oCKErqHEbw3GMWL/D5qKRCk5/A9YWzF6oQOq4EqxVx1HtO3CKf7R162/wWk4JR1LSwGVrb
P+ctuKA6WA6qEOidbRZCU9IQEBrZZOZWd4y5qoEGUzaOFmjHmtrbnnwviYgpTu4soyXLS+chO4we
KT0aELmcXJbg4lmXQVi3TnngXbfduHuZqcHvvxx+OS1je0RrKJlvJE4j+cVHiwmbKUyo5qOHYYwN
bJcI3ghswvZ/WKRWVwTNqKePA+lj4IK+6HfyQQg4+za+hkyU+0KNnob7kLeiDdro/pnE5x2fhXcx
4kPaawE8f4fHOBataZZtiLiPMOvSdYYV+kbhY0J//1idXnWPoiTEZahXS1OvEMA82WqgYvlA8xts
GERM0U+qJU3n+BzsRSSn1BYi3KRD2ZizqgBeTuGgZOVAQuxGMex4KGyGFSIMjK33Y8Y+zr3ua7+O
HIu9WyKGa4pfu4Gj4K/S28RL37zjMKl5DHwrMjbfmbUlICHDsXOzCHFnpYMDSL4b/rZaWiFldfPT
tJRh76HagL8uSDsu+nGNykbhsvWHXAjkdMBPRVp2i6TOBfcP6MBYOjERghjwwdsDXYKytxJ4FNO0
cq0QHhGlzZxVK/cHk5+5LDrme9NMzBd9IGa31eyo7Dnx3jkze0Pk5JiapoJsi8quca404nDqKWpC
4+RRPsxQYzGimN61a9lSmCwYft2iF9DGAG/X0KGvgn933cqMgpYNG5MGyZjpwGDpcAakl/8pei+1
XdgB8AqdvJxiJ1rZFYZd41ZSV8CMUYmxWbe5QX2fKg1wjdif8E4FrpmuiWkzMlgZvkj+V5NAUjwK
n6j404YYyT/S3rpKdZfJLkC5harBnQQZC9PtOqT+/Q+MXEA3s3xOeLweYpDhFqPsCw/zG9n3vP0D
Ohwel6CRTgBJ+A+zPJK/Whz6z8MDyLbbHKDmrfwnPpOJvDo9vGlTCKb8GVy2P+vngzFCLxWn3iP6
dzxw9rUzbjr9vsYByc+AdIHKCWWTi8c1mlksV2D/mwwgTvLy/hrXxUAxABMxAjb8JROTrQb+IZP4
X9yNV2SUfwVWPlmjbEkSErhjAQPaQqXbFeYpmMHvn29MzMevWr1W/n2NhmfMykHF0NbCfjlLnhf8
lWGsVrBCytHsrqNXFc9W7zZ8kWsUZRN8ZY2e7TjYW/z3CbzqAtCYCKJ/HZaxIkPQlSw6yFqsYVEx
P0kVVFmnDcz0m10rZ2Adf4FLRjBM4HaX0SAqFGHj5cb6WEVv1eHYBmIvUdm6PyPzmLsqc3jcqUwH
lps2DR86QGTitpmN2vmL+JCOkTVVggxt3Umc0c/Y7SBKSVfweNzl38WO3KDXfeSbDDc+P3Riohxu
ZIe23syeORWJ9nwfhkU4Ecbp04Fye7opapnPr6E08XkkVLlCtN2AQfdXS+zRa542L2zpE/wcSW9E
ZjJdIacdTDKRwGBjxrD2m7yLZNaWwAtgB2sMjBo1emboKMRwOn9gK0BmCOptAgAKKugNJBOnfbPd
2WuzUsVofUFnGb9aNAufo02EjbfR3AugVYWEM2xbYrPMFi3ZAu2x9+fo3zEyo0Qw5fr/Q9vDuZW6
fdT2J2azBvjW1JEN1IBUHWE3taQ9pHHTh0QjSOUcfSYnpj7sn/F+30E6W/vBzwinHTU2qbmi8n7s
2rnH1hAs6Q4r5xMSuUrn2qoeFIds16K6yZjqiL//F+hIFmPuQBAVe65PgaUFL5HWw4OJzg3I/jBI
DB2utWW+jTJaewgaNf1n988egiLy7jZCCTJHp7rhxqreWzoyY2t8b6sVhK86FHxaoLxEYyGgViv4
3bbgTv6UaiBIvsqi1+qB9DIzW2JdIZuIYb2TucAdx0UL38TZYGkZfb/vF5BOe8IGbI62XxywBvlk
D/9pWgc/8fMvDXUx0+YHsLY1pd93FdiIIGyS63CCEE3K/mhuiNRqik/YqaPcwzrxXNa3tiuLti1d
VVkGHSXINzQvXPJeM3ov2g3GnlKkiGzWdtFbmqmcEYYofVm08O9IMkP5zeqxwCd8Rhsd/Z/Awbw8
3zZ9MUPtDMzKRlbHa6+3nVk347NqMzPXpUIJag9VP1O5kytVLiWESW77IustSOwXCDSJS9x5PIfQ
+Q7FOq/6pnEviTDN2St47vcCD7iXNkXHGHHLODJzzKyARAoerR5JpK4nmYhcJL6sRAZ63DIJc0Wo
EYq9hfsaY3CZ5WaPCwjEmCdPKqxiGbbda9GOOKG53cOc5SFXGQtWSFufEfn5jV3+9b6LS69ta62Y
Cl2N1T5nkEVa/kJ1p6FjuqVlW9OE2LtM6E5+Y7JdEK5Uyj2AguHZ5dFtH5hsv6zw/ZVdD8esiSFZ
n5QjLPGfjElA1X2HFuT+xysmaBNzZUoZ+tc1O5tZXorBARBc6gPFZ97sH9P1KCVzSuK80wIQxDa2
8ImwfJ5oMl9a3p9AKkadnLuW7IHpQPyrDyJuwzAV4Dt9Dvn6twClJMp2S7nx63VYV38mwfmOyOmq
uffZEY0FsrYhrvhyrSDOF/UWd9DLkvj16oG8Mz6QgrcP3bqg/bEqW5UcVWpv5SeNSgubMAE0c/f+
5bnmYu9vmdcaqX6BGUbcr+Y3TcAQ+IQ/svyEVlRokTDVwnvK+bqbH8Y0/wECWm39FZOAC85/uBLf
86nSGPtzKZM9innBr1xuUxx/Svay+3R61HaAvBYyVIERSxozjDlJyirBZGVKITBU8lB4vPlSTEGY
9ZlApBz0rOi8ZIF4jiBh050/TYvL2bsQMxePacH5nIIxskibq1EYgFCUmwukM6uA71s1ce1PhK7r
T9+VPmOzZC4T/zKvdcPyyfbWjhVUQmNDty546lBx2tn88KcnlYMP3B5sdQixyARjtqtaBRkipQHw
KNqxZtjD4ulkl8wphYy7Q2DcbU8ATcQgwHfRrWeA6Su6+ariAPcLWV0G4kFUx68wsMo2m0h8IIPH
5r06pEXlXI4CQ/j4eJNybE4fAihxpvePXVHXyrrszzGhFUXotskQLfDPaY+vRA7Bz1criKbbuQh2
uAb4RRYzZq7F6XW0o5UUvQc7wWWbgujoFlwl+LlkMNTqE31MTI+0ZcgUV6DG3AIxsonutrMjGShy
diP1CfOTNCCapj4olzfqX12ant7XNx7PWfzbJrstlAtFyawV0eTr56GzO/JzP6uhvgblNTmwGkPg
UjJXDOQ93XIYIFQeQ2x+lSoy2a9iDGjgkl1pMBcYVEO3qe0YUsf5wyX++MwMQHm7fMRVODj59JVj
saLnlQh2lyndoW0bIT4C8YxfFiSgpIdM7uop1Dwj5PJcwLR5umMsYEtstyig+OCJG0Gb1WeqgysZ
IYcJSikNvJlFejH5ARo6HO8BKsgGOfZ+k9tgwR9b0E2dMNTcGTe4EWnFVw/zj4FMgfAm9esTD5mU
OTulQqJO3XJXhydKZN0xnE6VNvY46oEiAiNYo/Jn8h6+fLtI0V2ERKzfAozirFa5BkA5peRCdwUS
sUcp3VwU37roxVpfj5MXjsGxFjgFyxg/ucyq8SnsL+zXEmMKqu7zE70vCwkl5xg9sTdzfJTwFQ8W
2wy95riYgXufbsErj30pV2gLof/0sEXu5sOQCuKXTZDDPprTpgdaAOmGZAX2++e0+ih6zbrl7qcB
sQfZsV2cyAAAUbQVTVFYvfZwGzGNN08lqgdDuHt6bb/VcaURt1/vUpWuStRJQS+lp48Kn+UteV5d
arktlGQ9ufTM+SOks3+kkFH1ZjHZK6EcO2+Qca5yT3bTNIH5DcuKi4fIGB+ahb8y0VNoSY/zoe8n
qU0aLBsitUyOR5lrFyThY6I4bsxG6itaivNSEyipn0YeNRxQArlW5rxiB+Wk16V+4AwSyW8j/1Lu
qI30y96TTgHwkgIN6huFzp7v9A9U7QQvAzD+gaW8seKia0IFHNNElEpJtAfuwu5iJ//X1Vy+Oliw
BDuP8UaPyvzhJey8GaHs8D5K7rwvGtWTHMm15a/yXFn13m88fhWzvo58t1o/u3SslToI0Co7SD6I
RnzFouXouQWxEtRjISpnUxmlYuDITzH5sH8DT734H4VHc70mSu0JL6JyG8Gc9OGtneMufn7QSiNV
q68xmX9+O+A2F9ng3EivLe9InpOY3F+D4F0mtWmPgX1kq7FbW80MiC7eiWq4ElDDmKMSilcY1Eqg
dldWECY6OVzjfO3GIxzGfw1NBG24bmjOAYH4hNWeT+/eOPLGBxNeaCBwn9wTLooHv6OVb/u41sBC
aKbhxwngfHazqdIVWXzmfdJ0g1CsRDkcwp6JD+pgGw0ZbrIRO+mA+2GmCvo4Vi5nuyYRfZ8Ywkdu
rW0htuYnM5qZpgL8jhLmFCqio86yae+QjqKLimCK92EZ040SE2asi/uBmQsDgliz74qtjeryIf8K
vBg23jPouI48QF59ofko9WmQ9nHoieGLXq+M55uTfpZsZrjENJ4lNQ7haL5ROUsBSu6KCKHkdlRP
RZgFOVS4z3Jgn9LwUQqALRUU3/XVd8VJJWkh8+X6ZAJ/1KHVkVqxywBc0GHG6e/AeHbKOI1gI2Ce
nkLx4D7CDCCKMw/d1CbRSQDX7Ij53sy7/XViXhVp/dUCe+gUdAjl5kVUlgKqwOGQXou3v3vKP4Lf
m9AshsdnIY3mtzSRQMtsIObwI629eYpuj2j3xjKD8OdCMNc+uzFX+zEplaai6URGNvHIaVV3TjpN
uRlTY2/LXssX3Mi8b6kLp64EoNojlmmYvDl08kHNt1l57VsNG0xvLsv5YRjypWJ6ddX1x1yU8b9H
Yawok8iP1cKhB1qqNntUPFQ02tf6p1PJ2OpAXoaSULHYxtzeyi+/s59/dhux7v1GfCCxPzY5DwgA
2l3452BHej9lvNjWc9mGzfotjHygPqQk09/RTny3P6cX/OG9bjQBbC0r38FUAOB5L/fHkNNHvSoa
C8vQ6GXNFyBVfaXXOkGjFkDtL0CpP78UtCkqp7jphYKx5Lz2yzFC9EELLIGL5rki28Pb6zJg/OY6
z4d7W85poByIl54gCQ9DeEHKU7SPHq425/D6eNsv4PbVxac9gG+GBl6z7wPiRYPUE61z+rdFy5a+
R3YzuTxUHmiZ6ue6wp9L9D+s0KJ49MB8zG/M8Zpwf5TRIMa97LrOUSZuNWnfl4HeWvhGPBoBDC/l
35vVa4nvbjvdVdY3x7l9Pfzzghakyqztax+JKFV59SQ1mcTclpZOePqGRxZ7sRPVvjKkPN2xDN8o
qo/EdXyBLPb5jSd0C2NOQT4D7v95LbfzFdF7pvGRKf1iiMMWemBYlv4Nk8vjDsKb4BFSPJswS6mY
uR0Ujh0q0At04KWffJDLUJpZ2mTPDur6GXKCRY85Vukr02HD6NmB4wTC+U3sh29pISsqcutsSktt
blrzfZNIIiYJN63496BXfRWIeodJuN6s3qhxsL9j0x+gnDFP2uLAK9ksygBnYTVGog1f27VlWjUe
Tqf4+OioPpiXAixCuP4TPjQLBrcxBdL57znhc+FiHKcFxf3mGe0nSE9NpbCDvFkzg5SNRthW7u4L
0QNtU51uKOsocDyK2r9t54HyMVwQ+x3cIQGl+30wrR7W6krriY5JB+37OrAgtBnLeLVT4OZFfTYr
Lp4Hmqwq8On5CnDad8Y4VK2YmE1erXxXieO0yWscXVGxs48gApYWdPI0zLHKP5X4OTgGOgHKjbds
BJKW8HuZ61BHmIw/jO/x2lK7p32m3wqsO6N5AW5EQZm0U3OKVGLAOz8fYyGrFDcoXUPb+qTIpJk/
6L9elNXbxrZZ+p4D2S2/OpQ3ubhG+fb2YpMSDKdXP1zdpLxfvptYopkGWkB939xwcAXjK+YLkmk4
/oSU9SDomP7cUYAW7Rn+390uVRG5fwdag5brwO4c6407UxpWaWEBabI3poMl5o5hmD7qK/veCDuj
UsfcqoocZvcuPvqaqCIG+v2tmjs86MxHq4k6a21gKUZ/xgAqkqHViv5lnqpEEiiPboHPylJx/Xfo
B6ZtzinLJnoVkp2mrrOiTpKK1DGAtPTiAzUaqoD/Qr2hmrVyyUhXlJW6N2uK2pEs/G3LD5eSx9/D
FUo3XGFAg4oyl0efpp051lpH8mydb2QKeGpOrlkp2ONSCDnAiLGVlYkERmaBvhbq3B8lheCwZuFR
hF56UsOLUTRq6Crk3+E/fgRMyp4QpXHpyBztXXn2uDNlAzW0pAc0HzaI4aQW9a1EkDAtgBRyEDFV
2zRqvxpmBEXQWVCjhDUZv1Hr83kDssBnFOiH2T7Snhf0zEGS9QLPwPOoULTUcFyXu+2TokV0mzlx
sudwRavX6kxf8Q5CLGzJl5Q5gv+6TG4JPzPmn159nVhbBnnKgls34lZiTaoim0SHTjDD91jB6WFO
4VI+f1cgPDJELPlrAvt9QWLUCXfggxMv7Aaz2DSNhZBbpp+IwXbc4Fj7WJlRLdQbuhW0P1lTE2vh
pBVwwb/QFUb6Ri+TVT80PeRuvvzD5mvqgPWxnyg08QAU1bR/S+pGcC2HCOCkNg73gzTIdBa6S43e
KjpNEIxhXK2qVIyv5eGc9enKOqjtYKY4zrmTQE/bDEDMvcFFBA1Br7IUlXg/IM26fpyCjbNIjLYV
71F0XXn+Nh24mwO3fB5nWguWelX7Tk/i1kOJQnU2mVu9g6NRYuSffgJuUSH5o98Vak+R+DKBvtgM
8c47ImF1PQ7tV6UxuZq5Itcbi+UD9ngG/SqXqiTXWCHWB8cpCr6LwtWDeNCZF4LSsq7Fn4i0xeYa
ExA/n2MxQAgF9sq49JfNXLqayrgUfJ0TP92pWyZZydl6AnWMbH0UPTS/Ph4Szs6SQnvf40Yy0kRT
KMZnaC9pCKs2//BrDHRi5git/tnyklgLoZKouGbmINfpkTTr3MjUJj+wuyKQVO2YsKVqLLZuC1dj
CnDRkdu1BrP+SHS/AgWdrfKuFoS9p2VF2bEDJlLwLe+3piRCKuKlwH8PIFU3udtWm2Kg3sFXefRc
hghwvbJhpIB9Z4C2IIcDrHnicr/Y2xBnyxbKQPs7s9sx/96WCFX2SHVrHgtCWWOdA0ni/jnrqopY
1azqI6F/TmqZWylPR3iLGniL7LolS5eihat/1yKfu7OcQkwoTwKEjZVRTITqceXm7zxPEtCGQ1YS
mIE6nH1M9IxZatwIGwSThoJS4htwJxGr2WiOGIOHw0J/3fzy6jgI8N7TRuOfU8WZX+xc69asIGwh
svFGqQg/TaZDmKe+zpV286gqynlb/b/GtGE1NEDDg/FYQHPryNwzm+NUrujAOdEIJ3jBX7pZDzOe
Vx0FoilctIF8FU4jDT3GIgHmek5aNfqiRBBs8SzgG+MjVcN5NW9gJWsU9Gyp7/RFm5nFHvyb9ds2
6pgaT5J52MfYHJoqak7FsaPugIWlULxAOIDY1p+9hC8EIprQZ70m880jZH1wJoNa7iEvXhXVkbQ3
DnmiHkyoevNNcg3TRBXRLP0xgw520nrveMeSrlq3rtrKQHu0VEn6yo1UrBGoQOVntxRkuzCb1N1Q
mFnz1Rk8cY1iPIRyXIWP3rUu5Uo+A0qIsm9zqCUkiqB3oKLO+yavJ4sCGxIdcf2S/BtsImeOjktw
FF4sCm2MCE1gmnP6+7xvEkqFEsEcaYGA+UdDerSII+l9T7aNSOYrNdyTITQ6K5/W6dV+1b3+XZh1
UAIQicEmzADEAU6DWDwbduedmViBslmC10ndsbNV77/QRtOQQi+HOiIKOXWb16uXLEp2daAkbXOh
bMv7+ml9K1glHYOabOZmLs3bv30zZwkLMewj0bbKDWamsXSqlZ82oaPf3bszKNov5kFXbagdicSD
p2ZXKQP/GdKxd7pZcbwryqRVd1lBYExtC67N6cAjnNaP//Qa7Ztixbf7+O8jJzsPNd7ND18EZUEY
SGdYmBmxMU643TN5q9GvHhNtUX/qHU+X+7/E20wTTSnq5gKcrh6wUN81VxdVVy5wZQ9WBHurF86B
5SONu7rBMA9qab27HbjQ0JfHBCWuRJMDjEXDUMjTqqLtiWNQMeL3rbTipFML2e6piHxvKb7CZoY8
m6Oy1SZuKJ8qUjz75eDjuyAIIygGxSWcTdmheQz8qkXHA5udgwqXRRHeL+JY1JYmnF0upeFrak8Y
dfxdzGdx0lHSiPiqyT1dqDZL4dlgydVQ8W3USMULztjjqgL7Y6p0NOFTDvZuptBrc146EYVw1TDZ
mfn8qdCKa9H4Y8hA2U3NPKZkxuSYMe0ZfsIG2NH2lt5G68R6iDHT2srdaUdknLDxJ777celsTXaq
yBmSd8qwRjhs+ic4ix3IPRyol4I1SvPpGw9YGoh+EdOgNcAcJV7neGGB88c5vdcmhKvHqiPWeU7v
5Cl1N5A09NxiI0aI/Bm3Gs0btSFc+SKIwcpSxNdJmN/wfosxYI7BM/ZCymhHd534Xk9O9lCRSdGd
vciDELyBJOaH866g8x7no5dbHSeP0YaUOBajtZsYbELT0QR4yMJ7fhZ0b3HWI0h1KJN+rASf0RWW
O3sCRvs2Xt6NlQPecis2SD1LpvHhfdwQsweWU7shuipNzszXY84gCEh/jwlxQu5mYGEAV0yYM392
jeuLMSIqTMdJOZvxdqG0HNokQaSVWVSa7yYgZ43VhlNv+AUTi060S2dBTx5H1lqLWn2df618rOv1
3qhasn/iLh5SKM/OhoA2L3OwR8VM9RG1hVAFCj63REbhtxgxVTNf815Am+5R9ydKVJVqXsE49eY5
cmmevt3gXR59R4WDq18eolQaaoM8dTAbuZmyEVFg8dbCWL/W8+R+Zj9GiyXhH8wKfhphKW8sc78G
kgBu4z1eNk9xU4m05It8f8ymQ6/Okb296cFX/PuyhLUj6COPzgYn8mY6w5x5NfN+9chmoiTMJutS
W5KpP1RM/VzBu9vd31f96OsBZ6MpFjtAxT6b0yFz/0xtC2gxyR7je38v0Lwigm130/n02O64tgng
/farF2pDyej82hsUt1ckLhl46JluZgwL/4T7IWENTkefk/vsF4QpmtUpyaTkAx4hHX9Eqpku3BiD
WNC99GRr/WkF74bGJtz2khziWTA5Hx+AClpIiDDX0Qp548v2z/DTqV9K7lsT5y2h0IXnYELxEqjX
ZXG0PGob61Ap93MgEXAtrgkEYgsyta6XbzfR3tUBiv/r6v2MvLonRBd/5WB4UYkerwgQM8yGbJje
7rj0RXzp1ZYRU65DkzhZfRbsGcuCKjs9g12SN3zY5JijnWd+33a+t/n0SH7xxug2ioCVUBx2fvrf
3qIKdXWNqkhrWnl5GTTClHLAF5Om/NC/nfqNbc7fb7y7ZDAfgcJZWmR9aLbos/oLQSyAej3WkAsz
Q5KmYbafkKcf/IOUj4OJBY620203hCatmy2MNXoNjdo0dmWqsfXFKsgVHEEuc7GWXOLvN519rV3R
fsGo4nUVPFS9MeQ9HEOYp4DENnbfABI89Imu9B3ESiD/X0ujW23eRoyDBZI9mNr6hFqPCsuwSAgC
l4sedar89RYR9FgVlUwj0h3T1GTfLfy5/0ys14Nh/N866V9llC76GUuTlxka6rL1FAXyLTo/g/kJ
WMHR0YZr7Fun3v4P4oEOpI0I3YpKHzE109Rz/y3MmXnDwMXDZTWKfvWii1Z1/2WTl76fcuy6pFuq
vb+iFFYU2gv5S/eyldWFxQY1jB/sG2lmmyea5zgPc7u4gZL5i2rXPBlEYoRZoRBu+1+TLV8icmsl
PFRXBN720/dN8y8EgN0uP3lc6eIu6YOLF7jOtYoEEHDlgfQSyHo+b9GyQT5ho+p0cmRZNyFwpTiY
3Rbv2IvYbUpmMtK+4T2yW9LiMa+sxATw6qAz1VIr2tx7eB9Ocq0b8UoqrBJjY60kpXXtze3fDEVq
9e5Htaj117nove/EIZbrf/hFiT7QnVpui5Shbk7DWoPqMTPYqCMeBAZiaOzYZS1gtYAhXH1M1O5b
bYgzSiIXnpyE+ANB0ucbsWcdt/UDRDuP7/NSDWgPgK/eTKUi0JaPuXuZ8kUtw+f3Gd8r2+r3CtEC
NhG23AbGp+4thmUtgllzgcTK839vwgxFPabcgKENOurYHS3wTv/V5itHjnBCE1LRpAuXsYs5ZtXL
bJdRubl528gO24C46WGgUv+F2u/EO9CUXHyNfgojB9xWlkmY1fPFyRCpKxeKxIXmBtT60F3uwfIS
V3QBYPLRqZELeN8ZNSSydR1Yf8h0rqOJ2glw+J8tLtAQPcVPouJKaEyDwMmWWzgfauBie51gIh4F
013arfNqdV6hS90EjLzWLa33x9IWa9AMmOuEl2Ti2yy3pdY6PEmu2fUwUc6nxcSy+jycL6oiq+uW
+Wb7V8Km2CBmJ9GBuVYr0SvPf5V//xngTHcjyz0VHxtz+uFZu4AxqtdXbiBvNb21TQDCB10y+PNy
rm5AyoppESaKvr17Ygd2FRBtEqe9rB5SpTBi7hyfohJGhWEhKAEOO8Hwa414xvNWceegVU/ZFybt
SwoLRdRokeSE0XZBq7Sp2Wkr6ISYzUHSI6fYb+xp3DQIaNx0sPf32pfB8XLerxOzA7l8KJKkQ+R+
sAJCVZmq8NmtBM9n/LSU6PdgmY0MDqCyxOEWdldNVTE6ATag+Osj9QvqwVapZ63FAK7O54k2/tqI
Awmbfn+fFHediUUoelmh+Td+Tdnc0PCFhY/vfzW39016/I1Tt8j2Gv1WucAALEh60rBo1Co0pYra
h66K2NWZq7VFRMmsiicv80cD1kkYO5V63gcF8dktN8xcpt/oe053GNbdUcOONvlDfFyX4qLVVc2S
w+iOywIFJ8La9BcJSlSM6RQfofZzBWuimZNqCEr7QY3GoEwWxpImuSNXA4DjKpmJYhFHcpYTrRG3
d8+wroYugkAU8o9KcQcXZWWJ0Lyps7cbC70dpKW87HoHNBFaqjvnHw+UpO2Oc8WyYWRRCAF7zIZv
L5QF7JErhESAK9KjSRN/gervO5g9Q+GMPofYGjHq7z66Om9bZOI5E0Un8MsnGfzvkH7cAZFIs+zf
qF1ipiiRw0XbzWJlFnv6FAfz18MKMNL4ReVIke9YkMW/3VaxnA37THVws20tE9Rj8PvoV7jeuD9w
xp6t6dIIbFwuIVbiL4AgxvqPWzh42lQVUQLDSxnNYzQk3IEL0i6i8F/r2y4E0VhOi247jnKBMiek
3oa+L7uYUsCHWwc9639/GCHMvimxIkVAZnJVrWa5OMUirBIHhhrkHDmCAdqKdfkatBeIhKlX5Pil
X7pGIurhmWRPGq3Gzeg5mbct1FUrn5KzOQZeowUGSqcrzJZug9fZeyIG+Yvk2kXRPKJZmuucMQMq
wDS3sYnhIosndW10iLoPiLNs85FDQ7TdQe0OZa8hsE2oJWDp54eGLSjzdVSBzoidnn4kCzHbtdOV
LsaYjZI3Vo6B92AdNkARCO2egEUNUZUDCxic36qWIdQ+ejFl+YNXheUznBPjO+sB4Tm2laE77QoQ
+lBwcTasvopqx1kS+WrM3GIBQ6MB3+ZBqZ3aRy4EOoKe50kEZi6gpqgqbJhVrP6YuJhe+Giek4Sy
6ml2hoHfjSPxuxvYv4ov/EaS1A2Gx2DCNvwxBwYfa0CbCqDTiZAnOnQD/LgYvzsm4Fz4UvjBsVH/
MgW5C7uFgby0zro/A8jYXmNBbLXVX0RNEnBjVtyqAH/vXSa3QgVKYdBkYSlQ3NQQNO0hnG6DgohW
ZB2EfKL9UYFq3hY7v28G0PPeSGUYV/+ROg6krpleL43VM6bzwnJBId4hnNgFpOeX1WJmhajcNsbb
fJIfLfV++tc7VJ915v59jLZiM77s4sLhDeCOQb/88fH7c/xeJkCDkjXMFm9iYQo0aIQfjGBTj7Yo
TMX/Hi1w5pQ3jrDjHGuuQ7tAWhZES0z8c89T5PjJ5HbmKojw6SqqKc9iEz774PFQq9rm19gREMfR
kkf2fs81COkWRsRy4J6Oya6pCFdlq+oobnPI1VMSJqob9nip+d1ZJu2y+hCwzNkmRXyGy1CmhirW
M3q3gBS23+GJJFA+/kcqXN+fwcWucMZpI0mjEAoj/33aBZH5izEUbQ0RbtWo39oJkI1PaBGdiJFK
vrqQTT4d1ZlGwQ5Y8Ij+HZxDKsqwVTzg7A3eec0Ks/P58wCGJ6D5Jkw+5FQ0ddMolZTPxu/mqJFw
gH5WlnxWNz4CCUW6N6tj1NrT8rw2u2h0W1kiioZaDkq9tbY2vhhdEqaYwEG5n7h0CAegEjtOTEaT
Q5aO2mZoAs2cFVnAZ2TQg30Iz7te3yV1JfiW7pE+N2LSJSxGHz9U+2TkLSB6SYL4FKPsPGGI9AtI
8h1/MEh9xb4lZzNGp++c4t7c1kBaPdlUVNqJKoyWd6E7K/vefa+uEJAN9Sg9WsL3V+JMNs/sukjR
GIb3NhK468wfkzSmCcmhHsdNS65yTdXass3DJHiJnE4J68V++IrlcUJyXLm0b7dq4huNvN6rt1GI
Dz2Q6lMby2t2iwxGX8ZZAcNzCqi49+zLD5z0GpDD/0bt/75AcPiPja0Za6YdVhV1y3LvO9SWjpNu
XMBx/e9Ecq2czmO3GyYwz/aCKDeR0BiP9WY/OjRunt8ijY3Pb4L3CCBj5JMat38CLt0skcRbSSDw
klvMhXUYlYHIzbChUXsysbj9jm/MJ7vSpSpp3xqiySCXBMX7phVINLTc6Hhr1ikHWLQ0A8cklOZw
4IE2n1DLE6sgvUI40crQ0pO8uX0WhbmPmb7U7S+a2pvi2kir+8rP6hyUzTWOmDoOJuKfKqNNzeU+
IXXbB2GKbu5LmOGka0huIPSQZcUfaXzX0Ow7JalAoMLPH8D7A7zsSwBDzwi794nm4XECUvLQET7v
YipZLl0bmAt46gmVDLJE11w1hlSqSDOgecn3C/uRAd5XddZ9V2ITaZe0wcj1CE7oB3vwUK7TBhMe
d5cJTEdZDny9JHCBFHCmoSJz5ZOQA3i0mDUbd1oaAK2FQwIr0FdLv5lFC4NHcAuLQjutq/f/LMwG
EOvuGrJxGizCza+pYR8zDLdeKJ6Rg7jLOErGlVnVtzLNKmta0DnT9ANLTzI+NskvZnwy/xqQE9XV
CFQVpdMwo16OGQYMfY9S+pmVW2KwJDDz5FKpe4AEg5Wc7kuJ5EAwKxbv6glGKIN/ydG8GZ0oRemY
LnWQQ9ba82bXfdQOlgYcKW5vpHe920ZfzWTxdDo9Vmzq3e+ohA2QQTdvTMN3cjqXxpE56fuyZWGW
1DibWk5emV2EVXZBJoQ0UOFcwSMd2y3ShBtZMwmDjcdhfg+i/NekQ4cT7AHPGCtMF61Vadc1QXdN
SuwRmfnZ1boz5YiBb5FWd44GeGsbquHPxRZT9UdiBgFGJPzS91Hakplni6V+I8kcoaTcCfKKuIBy
AqhItzBu5XAKiBoDNPYpmkicxVfzIpDuJCbgEIuBGZqXjjjqfbBuAbgAqjpX2p+D00KetTIGizWD
Ps4Tr70sE/FXg2Oi6OBn9wZRIg29MLrbhEc2FmG8GgycrZYT9c2rePPFq6TdX+7cR1UnPmsKWbSr
f6zs6lGUHNXW1w57pfF5GzkIUWPr8qGVIs/6M7Y+RKuoSOpaxk29qL+TlsusN63TJhbpztcHfCg8
nh5mIL8ZpguBWU/bCgtGzQuc7c8gse8LOdnPxLCj1YU7G97tdXgL34eXvoFlmd+dpAppcuUi03Hk
+PT7QHB8pPy0+aRuVc8gESubySaBckvtwAmuDWfySyoWF8v6pm6MhO1JpnrOqmqw0LANWDlBrJ/3
J6pr/NkJirBmw6lfXtzZZowh0zaqK+o9w6ODcW6m66Ye1kiuP3wm7OhvOndGqhb0qAv/eP3GOmul
9GncRRhXMv3Oplq3dYDocAGVmHm6MXSjoYUOXgXQnitR90U1Or67oomqg0eGK04o3WgtTvBEep5j
a/HfUsBCH9xV97WWp/0bs/ycPE97Eq6g+iyRcEwM/SzvGqNT1PoGExGXKKREvjKEZqi5RTvrWnLX
AF8uqZk3y3coWY/J4rU94XSchPbmCoslIkVG+MmwxT3DPKhDNF02pvthgoI1ildCT0Ew777ty7HS
G5vWFCpy2ym1oL3cDhJaCvZbH2SH5Mg0X0SDS1HROSaBYLNnPsrb/IHeHbspXXzc2tR+4qujrPfC
4IBn7WyQh5bKZGayFKwia2c0dKmE93kLto7Nk3aOzvBbKf15a1IZeXCpT6a+cHohOoAcObKc8MnV
C3fMKXciwn/VmXPd5TCY58juvd6kq7TCzRQgKF7EmigI07m1Xk0SdAVIb9Wkd9IINxur248lLLHh
mf25Zf8D0IWy2/mxB2fEDfJnx+gjKNyyZOpFctVgl14NAWG4s6JN9TFG/f7CMa0YxnH9icjzEZRa
3HoedVnnVT0AFDCJXiagCLJ4L6icgWR51X1iW91VH551hL6nq1BKH8L+kzpPMDvNXxih1d+Lo+Nu
USiSj9NtOGMwY0npKBYyf0G5tWt3zVI6YGVqcTEDXY6V+XYtX0uovjxQ1ff53qXDPSFGlnuTdWuY
oqywZWh8qU1vo8DQxKAFF43dOflMf6f3vQmy65n4UDi77HLqRY7xYz6QY+N8PcUJcxGsNbkK5LLg
c2noacdguzJyUxyGBF3VkMI0+syBiPL+w0IhZkoLu005FzN0k1BjWAudCipTQe/cXdw+paEcph71
3ZJ0avuKQGYy2IsOe1T1s2P7yxWzAq9sP8DYWkGtb9Gu5/G4DXxjXS4AVt1QqldohdEjLiQlzYqv
cAgON33+hNtMLWV8LWb4sMMDLDNv6OrZPaWVCNx8he7GQ1K1BKHsG3A3GsEbmn5nhEwPY8M4hl4R
0rZJlu6rQAInptqz5y9++N1mcx7BzqBe4EW+ptkB/dNAlYYmSwMQGJ0cz91um/F/9kQrcPLhrywt
lQAJwMPArr7H2cKId6gCEWfSOMUh1dogbhhwW6TGsnUCxUQX9xz+nujGQt0BRYutrCftjMWdQSGE
/DwxdQcQjrE7FR3VdBczV9qf0JAiFQnHQNPYt46Ib0aqeNEHHd4p/nurqwKojkrmOmXSyJtayC4M
/gHfCt2oyY/FTTPB9ABWCUbriyqgT5u9rJ6H08DQfyy7S/tEeSPqL5uyUOqxs41bE2ZAID2kZZkk
HhP9NeJh5Mkr6cefZK2NlrlNXQzPGgFx3KitgoS62N6E8k8fkitl6fUPy2kJk5eOn5szCzrOXK2w
33yMdkbnWJRg4u/11N5toIc4/xKDraMk155NarMcKizX7wBRYBHfxjOPDBv00VkGDd95JL+QvuCg
DhCuX5N5vt7rv/0rwWpYJEA/k/7oSnDUVGEd7JWBjHH4QdpfFiXODJAACGz2pwc10FzMKUFykB+G
q1KAuXA/zFdkj1+ZsLOe2tMAUFrMQCNz7eT1yCrUI3/RUxP4KCnrsHNjtU26uDf6tOJiZc7cadH2
q1neCsISlbUYGwLY4tlfv3Q/V+ecDWROiaxOIuxK4GhVmMu7iyKvnKwQ7IFQTRRrKdMm7I0nEL/M
9YhdaRRQr8xrgnJ6CKVXRg0XJMI7HlguVqqopUisTFrHumQ4vqDYFviGkL9KL1RUyQuQvNNyKhz5
SPF+4HkCJzifwEqTMxRZGyLQtLHKGCv6d9CQSqLpgslVnPeG6rtJbl0gv3i1li9tuop6QeMvA67a
EXgaGu/BoMHhMQd7nyC8xG4m8CQkCCwr/dhhUmtO6zXqs0Ql9BpoNuxM47402BbzysVaTGTbwZew
Db8AirLEKi7MKRBT+8vHcPUbk2fBOgMI9mw8U4zcbzpbS0P355ePNO+2dB69uAox0ozsjWtajXAO
SIcZUUs7oqZOO+MbhbtGSo6QDBPx1hwoVEF1mfW7AGr1iHny/Ujnq000D4XAyd4vAWARRG4sKvlr
jPRZZmyciI+SoYdIp7Y43pklzb1OmGooJp4HpYcBCMhD5frABjoyD63Z5lNt/zKN+iZTnSTW09AS
5O4v0PYm03KFubBMJf/5jv7jNMtNZXavHfhqNmbdKQ8mM+W0eBOjadlbY20OyfFvHOHec+eEG2Zh
hMP6x1MqyHMIAgVf8d6e6NSiSTB7o61wstuc59nqw8wMaP7M+gsHellMGEK5R0kUbh4BBnmzhJWc
/yE5lOO3Zzzu+fpIyU181iTXJgCKXlmvjZ79Ww6AN5Q3OnYEZvHdU82CVE7gulNsKqOdDkTcOdNG
O+q85kWlNgrWgevCHEH4DZJVe/D2c8Xlom6D6EqptBWNe4sEsyLaP7mRLCNiNjx4Ns3ZfWah62gO
wu1ObEewwvpEK8u3ZK/MiA1+VFMNpLHAHT/qAsFsra3a1GJndJIrhP44ZSprZi3OqfuYlQ4ccJJg
LbXyog5CcRL3410UV1P/13g5QWvm5s+yo2DVMkv3WMuDPcQ3VXFDDpbWjf7PYlBfEoOMOAlBvuDf
BS1xd5W+o52uNp4b30tQav68kEQMs8WhPRpp7D6OzCHpe4mvIWt8bi8qWzivTS7FG5b7HgwW+YiE
oYd/V0EO02amSNB1kA6xQrzcy86SU/MIUV6A4XZYoFpWuLTKaUNcRtBm8S129dNUmZ7fHQuWlW2T
+71s3FZqESckEnz3LyP9/l7/VCkt2Z1SWt+qo7wzxb6g58qqfhthPCcFPLSGOE2JKVjWK+p2x5Vv
jf+JU62hYiM+7YRGlVazQRWsN5wHgF79enReMfi/EbjV7VKytBuoEwErTMtMhb2DIfWT+b0qOaef
4wHNCpFkB7elvDdTVgAmoqI8yIfYrD7Vl4Hx5juNyVZMCYPH5sfVhLCROs+Yv/Nj90EDy7t2X+ue
qCJ8kRC9QLC4k5LLKYntPvJPRlkftyCN/Fp6ouiuhOzu/OrSVA2T52tcQD44UN4WwH/+h5+COwG5
mL+/dhoktP1utb57XKpCrG1JwHX5vffDAofhJrE9rOE/Mj+3moWBELBtxOAj3wLr1PFSMMxvFXx6
gDCdKbx3NkezWyP/Gl+kDyrQuLmq5OY34Qgy88YQKKDmTEYee+C3J62cLaXVEJL8RtckiSmO2v75
eykUd2vUWSaRPiisQKo2Ovf0NsFDVTsEh/jaxE8+RtNf+kq9QKb8EguiE8dxq0zZOQbIKWa/LeDs
qANCTso1icFm3VE2yB/A6J8G85Q+OS55vjTJZfK8uHeqo51f4rAQMZuwO/hB+9ZWDVvHL13h+pHA
kTFzbNXjwc2Vq0eZH44vUKl2BNJI60Zm7SzsBQt4ohRuUEzSRFNT6F8MEtm/T5k6ExAYluDXTwyE
kEyqmfu/gQNXtXYhNUJaXUrDxZrB03DoOnAs5LRKVlwAuUzkx82DcfMlDtyIDpx7Jgbupv0oWVXC
XawqsUF9DiWXjawSiLD3QuQz0kCbYlGNw8hQbh637kwK8Q71s76xGny5s49pqLb6Di38UhNTdbzZ
vMvolkdHsUq1xNLTPSJW1Wi9VmJT61+Ka3HP9aoES1VGBgT+RFZtcs6en6C96bpfo3iS6VzdWw9H
YR+oT6rQzoMXmNrQ6P7WVi6cFxBYHT1J88jiO4g15YypSoUY1n9IZYSn9ApATeivi4qtajbhKwRp
IJKB1Q6fW6+n4mj6iLqioe+XgFhyqfN1cZsb36yB5bj6IrBFcf0Rn9fYgh0u93Am4OQlvlP3T5in
JvGyRFm4UXg5jKXkS1DTp/tKc07UR/0ZV/t5hB6S/3b2WkIGtVCYFmxRAiMLL3DjcUt0kaQ7M9zp
98f22Tfxf2fegtk7oCd2vpKHo6qXHXVUCKUZ/27SuupUTDz0eGgXWjtccEsgCnl/8bvSu6KpGBJE
Ptav8DDG0PJFktZfTwtd1jNu3UFWu60XwDAMDgdxdP7JzOgSc6WAny3hVD37vaKTwFSsdUpqwoDH
tfQt4K4Jq70gvcIgnThm7r38nG4di7IDjYacjI93aZyAO8xcUwZgdhgF7BYmrZ/a4Zw7qzx7I0R6
jT3i0fA09vVBLbJjjQsNIurvA7sbJNEcykcnfb4KUYgujXzmTiYjej+8DMigig51r92xS2a9U+Tu
0gCGyARmm+eiykeZi4Oq9e/97TPNGb140eXXfciomfdlWwjJr8XlvRc5IKMxyZyX2j8RAdnJQffD
JGkFVYU6vvnfI4VN6pcaGminZUbWIgGuGxCr8UVfCtpvnoF7yOjGpUFvLqOnvr1vVjCaH6aH7DV7
jNWyUocQUth+6qGUmnxZBWDayb5dgz2r1sWj50QiopGMr9MQQCmAJojK3yeVhnhE5JWqXdT18IDi
cC2drpLnUqJildEHi4CF1Xy42DpBh8fZES2xhTb6OmFdQJp/J1cVAi0Da/7aVj9ybQPqAhhfnVID
GcWyNIgMUtAxMvTGlw92LWE2+Sn8VDKwbFuAZjmEEpy1j9r4BHZTgWqYzO0kaj4XYshkPFP8cOow
L0OL7prPrNq+diPWbnRt1ATXFJVFm4EnLurjb2LVaWGH5JV94EoxPcq19Z9k9BzEjtnA06DbP0oa
ICtMYJO5JZfUO95/SDa1cQC2r9dV55ukV5tgAIERhB+GjWkeqPVHvCrYjegKv0aOh2ycTOuNMdYL
aCkAfamIzuEB03w0orEzD6AMvZjDGYmlaniqVeHyPjpCt3yCgYFNUTQiwcZRdgkg7lL8VggXKuYF
r5M6W9BawaLLNjFAwT/Ba7RXmVKL6HaFrxY6tuB5+IWZ2fBv6jMQP2wNTAO2lkiwK2XygqJgQsMI
QwUN0QZxWgzlCj/PvB4NUo1t/6HvPXhj705lv5/BCPDAVygPO2x7V6gUnqn43Y7UprjwoAf8yAqR
gxcUi90Zv59uit9Rll1VL+TreCseqaQjDrxKYLgYrz5cdCPy9lzWpBuL0tFiXzymbVrb5jRr2tYy
2RtWy+5pNkx78ITiYJcejiO/9H/MD9D6XN1PUbS/kaOySTO23ZuC+DgmxfpQkelN94XdeDBNfwiB
DdRK+D9hxH6iP6H1vJJU3UTWTgz3xuF4qEpFaJWLxAPExpDAvnBI2+EFv2g3uu/FjCdFPNs1qg1x
3hP2gQMHOpiGs+M/Wq6ZpiwK1FRz34aht4zqBiRTrhYAMBCYpU5kIAUS100U4lrpgTNMyAw9radK
d7sPAMr5ZMROOUijQG9658pTVJLUnDlV3Z4ii8XJRvbG5Ub0SLf5auNKxypKpXgCBR4QXvYoFcGv
F/NsK0mIfSm7BxuE3xrgsI98AutsClGepX20/+9wSHqMQZQ+qRUEWeTtMFppqAeiwWaMf2nZ7L3j
p3/NQmLhDk1bnYXDlkNETerVvRnGWjxMvykrCFLF0IypLP47EaxTORTyM271n8U0NQFJh1jwmFQx
sOYJYvRC3DGUoGRsfE4RUwbDRPFiy7eQYj++vsdyOgEgiJDEWBjGIzackYR7RU85M12FYrI0gZrW
hL/ss3j0up9wS46kYVdX+Un6BoxityasMIuqXO9eRBx4mPXKAJRg9hhoIdGm8uY0ECXLAUhY772N
A8LRbmtWVzndYDLlUR5WRdeiZCyd4BK5JPublpKglHDkBzGgKtbKZMgkaW2wrv/xX2hUeGMxicvl
iKk6O4OEVeOJWuOSxxV5bHfmvZ4xrdm/Nqs75CgSzQK9YYP/jqa0axIJrdNNzf8fqoY1oHwMG5YI
+3I4Jjn8IfP//3y1LPLtcGH7RiOa8qmH/kZ4BK4obHraUtznwsnvYXMEb/yFypoisrqkgY8dYp1d
O27/gZMgTUYSpTlqi54tMyn7UUmD9KEmq/OyEbMfkK8uqjqacoJIyDakqkBhqJU60gclt3PWOvt2
/h8dZS5DnDNpLsXITF1vb718yxI9UtUn9uVKgu6BufbHy25y3vWP+sCCfpM5Y3KSp/afCEbx1dwa
Bd0P9FQV1kC4tepAu+Bwprdzd4ovveNZIkBjINiOfFgWdWvww+pln17YBWYzUGXWEYHw+2nYy1sA
JlSRwjPpgZ58tzjgPuOUk4YD+w1eQBv+sjvQmXILnA/qpdS1G393UFpBBn0GTsNOWsbVUoxUn97o
zXcQ9XAToFr2tyQXbrHQqiXBKWSLpulXDENLItGcWMJxHtQdiWdKlEQG5x8eF6vSZh3bWPOU86c4
B0t0D+wodXVnX75mYtEirq4htCQYhKR93Wa+xUJBUHGL5PeFV89ooV6QABnSbFHXByJF/dJ//KbY
XeJV0qV+iVLtjiqraSxv5vYWE5pI1zBq8tQ9IOGDsx8oVkQeSx0efJsCfbGMH663Xwfcb0XTSnzi
Tov267Ng6nu3jSFz+9WoKLQUdOf0j9jpwVWxAEMPdr9UiRIEfm2LAHDJJ8ZoQi9rhZk57mRwdh/D
5RZ06szPsSQBTgVV6HWSmadGo2Lqp5UJGiqAvLmt97pjFtZ7pvru647yORnXx0i0gBrkM/TLaN9i
7lWFJKpZTLC+U4nyhyyRZoIzwAmZCbwAzCai2OvVqCh0iOmLPm64YImlbU8DIl0CylPZiTmV5Ura
o+2M7jio9gagtHgmaAiMCBphQrtscF8dfZk0TRP/iY0Ng5tegx0HlJPABV0Ksu9u4022NIe42vIE
fRMF4nnTfnhEbn9K4A8Cf6ImnNKpana42enqKBwq9NoLcXcOxeNJQ6F8Uc5VpCRK2dyhA/NyI1nn
lypnW14JBUsIcNbwehDRXgefa0lXjHmaVGwEPrx50bpuNVukRpHFl0IM27b5PmMTkphB9lNts5Am
4YREcxGQbiv/dtmzHttyYc/xPrHLg67MmCSaLPayB10Yro2rSWftjBRwhKYx2OxbPaVV1qgS0epl
AhJX4R0ZE0StmWlBGLK0oDz7q4yDJ2YmgTlrB8GAVzcHfJzSdrBO2ZED1w3eT0vyQcT0QvxGlciK
f5oeMgobLM2USq97nfgipkypilrvNw8Dot8IMwsGEqnKjRhFORSM1qsMgJvRbZe5+2+jnBQXlBMq
pVpQu1moqZ9Cm2TI49vWBb20psJr1tPLPUGtaErkX5LL1YzwIj+fQlF176TRPv+BnER8Y2uhh8LH
aCU0j80SrHZDJsvZlqnhuasFPOQZCeXyp0fleMML6phLK4lg0pEDtUF3MLkgqZKH863uVzCoV+Qm
V/jpF/U8Qb4E/7lwJeB2jwqZ01OpaqAQsXnyLU6lK2XtGFRQE5qtzLjsjpuYN5SW0O4mP9z3cCzQ
OOOat3AVBTNjQcrlfjrmUt1tyD6cSvKkI9e6By0BPqjo/bv/0xFA95stez1/fb5z5Qig/aXzI4GP
P+Io9QaEtNpOc0a9pmbBRNrA6SRIB+IYt75ATIki9b9+rqhAGBSVRFydwBpZpgBkANxYcrqPcIcH
VVxM+dVsGJzN9MDNIMYjkTdm/9VxVIaXHo71YNENpyUyRUNi7eazZxZnoCVkKPxfxoiDWqRr3vm7
9UrmtGWv1QijkTvk6fqo851ok2GVknDS6oi2ySvNpUrR5BI8pkfdVGsjWHfpQ0vU0qhScAg9fXR5
JdmcZ6G0hdvSpmVQ6JCEDzQg4OqBGi6MhLhZuwmhNb2Eb6Tf0iWwVkej2hz8NT7wcQJtvBWHBVCg
r64JP2km/t3B3pZZEl10E1PaMn8XFBT0p9/IwFQl5rDhXvpjAK4xobrNykzPyZjVHx1oNZVfHe1j
ZV4q+GRRuPvpXsIivk39V8OJLZeWeft2E27bvmKfzfEeADbT16hDKMVH9lK3zF5ANhxxBkbtWxau
WHpuGULVzZAGmlpiIPYYpntu2MureBYKKsQju6Vc8gsL4bdxk0xFpSNOqFU2BYkb+RXTqm52wI8d
OtNLVtL1PR0ftbhVNXj11l/frhZKXsb5vxW7p8PzFTL7qgBHjXakRf6gaiuT2p28MkBlOIIiuuzf
4w+t1tCTPtgruEccT/UEZvl9qBjXVxgSXr+tE0Fqfa4uoIUOPbbWm6AMSlagQRzDFEhFGowzyFUF
+C+C9BBzi+yNIzw62MLRALX0KztrnxSUiph7sJ3t7BwwxKurCI8ep1dciyOWI6urhBJHtZ+KNpUp
R974I98PX0+KvfjisQGF/OzyEWv/JcDQSZgHWfNazJ9UDHWDkE1tWXmxLc1BcX7pQk8HXwDAygwK
jRFmo58YrkJE24tQ5uQlgSHFsXeKImaewvAyYKKCDB+0D6uF/Ji8whrlrJQeOg7jF/n2gd4haztX
DqOQIjyp7kFee4S0rFA0IaljgN3Anp+N9wsbconsRu4Da1roAaprfAtD8GAzi3Uvwf0wiltwEDg8
nccUtdaROpVfoykJQfC3Xda2nJjacVEMYbBha8nSpNYCSmfIU5/tNFKwd6kWoZ+RJzRlXRRmwYgb
IxyMXgb5Yi2vatSUMKBgTpA+4uahzxCnipTHPg3SzdwlYM4UWt0xJhbHg/vCcLmAjrx5vJ40qrZr
ASW0x6Jrub1cyeEzGPpOUqkVRa1jf2BKU9CJr09waxsvU9e1J+iKYhcFjsfV37NlJjJ/bUNp/R5K
Enlj8TLT2jN+zt4Odq7sjj3emeLfBNldeWKf9l+Ie4qYRuHyu7CLWVWmSPuoK0KdZAImhvKBwBQk
M8uK7kKxdNcRmQvGkyOsPj+sa/APB47O1QjvayZK4PVtNn++bC+oUm+zH1m9EJnU3Uhg1s4RqlT/
m62ngyBPBFudlXFdIQ4PbyKubutA5JdoG9vEBp3COJQ+jMCC4s59vD9yXomoKKtyYxv5u5/TA2Zc
r+wcUOyYeVe2RFc/tS+elzz/TwLBf3JuIsIHR4pmHp6s9BUKN2C8jDYEd4NOj0ejtokcOnJ/cKzn
TictHuoyZ/vRld70GtNS7oVPXJgKw/0m+X4FYxkvYdwA21Ja8rSzy8S1XtyaQdNlHnGIZlgtVvLP
m9HLEo3Sc7F0PWlr60M03EKWeKuvj9+QcVW8vus/EN7LGdwRB6v0Z61Ys7ENQuGkLSBHrjIywWlU
jcYTLAXJeJR2cV8MboYPELyD6WsAo+r6WnG6XGLdypEJqyqlQ815lA/KHZtTdb9dFzSZHQqUQcHk
Mnczsn3MGfDKoUHLYDpMb9w4vgHlP9qEW1nhNp5dHxD4uz4jOnPn1PcRX2SDszGGKUS/hbpTM6jG
IqsaWr+dvRubpw5koZD7Ecl1ip4UEAf4BT1UkDxzo4hNphRqufRkauKcorGtAj4/tc2kpvQMkf/l
t9lnZ7JqmCuS7bdc+ZGZ6xZ/QxHHT34sx76bB4iv1kBXGHGzBErXPbUC6vOKLK075s0LRDX7AOl1
RyeoGotmUJjknYDZwbD59HqGSGU9VFIQsO3O3FXNRXCHSkowwyqJs7cN4teSsg0J2w+UoPFhwF8x
UFFnsvte7/brtILh/oWaFRfDmKk2Mr7QfbpWAEGhm6uABVDtABzeuEr48ygTH3UfEE9v4LW9tgbB
caxGcl0cm0FXZ7V/+LgsWMJ67cYZif9dUkbsOKnIiDekJL2GyWAtcArlY6UPU38xoOjIjTSTykRH
iCor2b1otxSeNCsPZ2AJZhLzTTS+WMOxy80cLzR202bcJMcY0DEvOPnVg+BejBTL4vIyO5j8AEg7
FMHqympTO2+RuMEDclOektaG63ISO80QwGVG4F/89MTZ3BIty4LRVbjX4KJyYWoRY436hooLlaAM
Hxn32ggho8c/L/o7Mh5zz/+2RVHoqoODn2DBaR118XQ61ZiaxiQMJN9VWfKvWBtBlFJTG+qNpytv
UguHqH1wSLuac/WNnpLqMeddV36ueTkXdQr+JEWJnHh591fwcMejoxips+A9mRPxlQeDT1vROTEK
tqKQi5v7XwFEYbiWZmQXMEDMXwAzc4D6Isszg2LYRt0mPGsBiJarCI39LmdhZCD/0kRKXWuDiVVz
dSwDCvNWSezqnfxHo+jn1I/X5VjPvsMWPjcTC9SSIpN8H7ax60iZs86uptMofGL8kUeOl3QVhnpt
zUdHcJhD8xCoqeNfDgTxlqqZD2+TSD9ef0+3p4eCT1FmUxvRRYzUjriHAGTrCHR3yGe8k2mqjlzj
Ef2OB1jYNnoP8fqUpnIM8aZ4cvgFti9sCp10Ju9xIDc0hLOzFY6yIaK60oZ8ZPYtlrnCiNLD7IEc
eBKUbU0qYpMJwAYlkPl1LnReqRHQ51WIfhdvJiC9PG4871HL11d1JXDPHEVQ4pJQGg0IW0jajl8+
ssIrRbs+bmDwwpqxtDmjoXkHdSQ52nBzWGr1KqnNU/0zr5WpbIkfADeKlKkneDJRPLcvKBrocvlf
X7in2VuZP1698pU9JbQ4oCBsaN/sOwmIXgJfBhohEi2rk1l/giYTbvmWKA2fzLK9J2ekrOEvGEIb
N1m69qwR9L3R0g1HRYExnmNRFlReDyyGeSu7qI4xJDURIdd7bAcFi06RgrpagogU64TOqTR0fhJC
C/ZFIFhAHKEFfEijYM9yxBUW2qwtc1dNfaI6tNAOrXV5+tQP9K0PXNi1N1uCWUMzgRIYa8mKvOVa
DunM9Cg8l8S4nZn0y3bXN3P1Km4hM/8J95BLP0JHbYB3QivExu1KJ3veMQhw+4hxfd4P2TTN9/Nc
oRezeya4qxO3N4Bxn0aCzH4Lp+15d3H3w0csIbQ3GPOZkS3qMWcJkC8Cq2gxaMMp203aLEfkC3vp
tR16iKlb5MLdzM+eqftNOg0dllHRkedot6c3mUFP7u4iUm3X3CHvDSr3WP+WV0voCGk5666Xw9p/
6tyTKQqps4WPgiiWNNKWciSzzdS20fM438Y79PErDsWx/28Zhecggs32xzDXwDT7CkRRaJ4IQaOQ
ih2I0fGC7ehAIJMDwWrPuy85E9mMg+3btl7e+xZPC0ZMEXPlLv7+v5eMmEx7BO87R5P0J601XXdU
Z5MsGnm+62p4T56dNFmdUj3qm233SRfteGm+OM7E5hGLYGMz9YrPRimwUDCXeRAGoowcSHp8vRCL
UMoaRDdG8dzE6yzH1sPscYtZVnEpW+HmrspVco0JmC0Gt7wRNMBGUl0q3jL8SKqsNTBSjhWCieLZ
q9+4G1im6ga+JF9GAuVJE1J2xx+03J+WCeqeTPbCYtb+W3oOskz4GbY3bf7dBycK6D6q6PHzBllb
mxTCGUDDut09upcVc8a/RIua4d22iq6yZbH2Tig23QJyCOLoY93ca2m+jPPGS0ZI/v/TKKu9x7MM
p6nHSOwFN5kCfSEm+BleCFd3hRam9BC3GbhxNC77gprqCyI1aorwc4iHescvOUw8t5IKZALf/2Jy
NQ3saMvlWBo7Dt97DvIU8EQk1Pqzz2oHYzTP4g3t1NcADdDV3/iloc4Cz2QaNL+Arg7LkcCbDjEJ
25dbzAkRrFmYKGLcMKjfbx6Pyrsf53czNBWv2xCXxcvuZFYvET7a0BPa4n42IQv/BfZKRADRwiiF
qcVPobgc14wL8pHMN3AiMb33FfbGTPpbW+ieK7E/w2vOknwWWS04qw3NkOHwWcN3OMp/XtHx+R49
5f+NsUqQCcxqjUzgGHnFm6t0/i5N4/FhdpgoAGAXf/uQW/5g73nz2/Smwt8851issi8bGcVYw0Y9
2VnMYgGjADls1TQVT5KoPrrPfxY69dVuP7tkDbZSSVWkQtu3G8TMxCDc530Cep0/wkKZoJ+wH1eq
bEqyhGGRB5J6xG4smIzV3X5OQy8HCrLiIvHQBRAKky1rBR+cYJXDk/VAMBGC1RL/fvd8R3qlomM3
gMsf/WWpfY4UEqxfWAav5ojS7V0wipLHFYCXCLTgl4kbLVJRrPo7asLUcfcX0AAaKhdKqy1tYP7S
SW/tH6uwG1R/g3lqITJ/aalCqN2OocpQ5ldg7/WqaSQrOp6IKgSujCMQzvvBlborLSixJL74B8SD
qMrqJCRPrtuBBCAQYpPL16t2QHat8hJtxlhjdOudW98KSUXZu/BazowS8zTds9nVX30RaVy6ue+H
lCLKOi3UHjRzGRxZ+/LtEQaf9aJmD9Ez5uSG8gjagcvDmgf7vgQJ9d+serK67wbsR90KWXdnoZir
qE85NUcq03g0jNbPQg7EqD98qlGHEneL651OCSZT1kMRAxUFRz0pvzBAJjpf5mbVCVR7r8NNYlRC
YcNkNC5YEssrhsFBBsFFoff/Z+iZNDu8wYCHEfyoKX+EHnNwwzs9lpownEF9NWzHUHI/1wGwyXIs
aMttB6rRlECMS5baGPoUhUwmDsk4jzgCNxAtoFQGVdMuEDhZzoTEw5pBzOhrbOx2ean2Vc8Tw8rW
yFRJ/5p76Vy61dJ/janNppr6tGdxocwk+TEZdeO2NnCFXB7lWLvb1TVBgTrUrkM98v5fVeK3X7zx
OTlVQ+5zO+GDk6HxiJwGycFeI3F+VOnjiYCx1oDZ1846/RGgBFu7pf/rtf3Tbc3HljvoJrciXJXc
fm7TdzN+fZHlvWi8L8r9HMQ3mdZb/AxxeUTGB3zF0DPeaHKE0fhFh7R+6vgAwWzRBPHs/qXC5wlv
DaEnz36irdUsaG8doM6UHp8Rgz+AreDApGwpSAqKsb/goDgiYc/tbpQ7KKKqDP6dEYcEnTGfpgL/
iJQbGAtFr394IZ14tUJ5w2ROvd60WX2xF/j/IzJHA+5rpj3uu8oA9MOqpDb/mxsap4FGQDSxblld
91z46Vbs5zftXsSVpJyO7SgKGjuRpT+7Cwkcn7oDjMv++/DbC5O5COh934lvJCP/uxwA/6mq208I
WtkaM1w6aWSFd5HrKQejS/bafVzewn8CNlN3bO0GRMSzisEl67zLnjXRhngbSYbeSZ0wz5EnvSZv
BH22Ph74zrtGTQD/QS2bmG7DlVTpoC9VO4FVtNwJytyrj6us318tWNtnHn/x/VcpMo8VSAr5g2RW
ltzs1KQVjIZ+V7WddV2XaJkgMOcW7ganyuohztuZWVxm68QdHtdtBfeA1RaZMEW+iYq22I5rd3V8
9ZXiYrTU/bKWtyTWNY9VPYlaWL+XElj4Otp3JCxYviP0A6unVnSyA/aorss+3nHzpwqhjC1CZ2t7
UyreMQ9o6tZZMyZMYPpLp+FayW5bNOE47XfGQNoYRILspNEC/HvrRWJ0XCCpVVn5sWdKmtakM9gX
778y492spLzyQp4DT91PTs2OpXtx77oGHWll7FInN5r0IGIbBCrP7+PSaeafZ+FwoB0Y8SAqL0X+
GW3BzxBWs/duy4SkyH7ZaS3Gj/N1uL5KuStn9W2L8v3DHN3Ftn1GkhnOM17ku5I9IUOnHEX4W+9w
fISBVx3I2E3aa7B+5qwBmKlM4buCX2GDmJoK54AJtaTSTRUUfA4RghJFMwTQsexrsxze6sgqOo+0
n48N8Lw559Gi0e9ichEbAYVaSbWKYzXNiyatzouopSsjaIXOkpguZhDIPFW3tkEF/iSo3uqb7cWc
Yb0tuDLQ1NFn+nNZPDJ1wBgmHC2yKROJEGayVZm0hbYtP3cTeWK7KX7SNHzorhpEWM8ZjBmgBTpK
ExWGr6EzgExNv6aRAs67uZZi418H96qgHb+1ADSStw46s3ipbdTGcT36OMjfBYyIbF+wUflyqkLA
NpS6Fxl+t2VMJPxsM5sSwYGJU3ugiAzEsiCZINFPEsbRKdw22v4N7rNpBdXE1bnnDanNrhjnzB5k
jW/c6pyjy7NLRFECBT3FXhEfk+W1LVeDpIluLqLL/Bbs8vt1N5obn77sGhSpKPVDQGL2VkXVPtLc
FMGChs3JcFcyqP1CQdgczBHOB8Z/NjReZRhHHlnU9q7EHNqkTtW0jxHkYkuUQMy98tTuOKaP8xbj
qZ2+ZOkH6IXlVgGU0yNtllaVNVs6uZyb26k7QPntSgcBRb0iPz3H07CuANXX5TxShnRxmYz5im2N
7+mZU2bXHtVRGyZGhmsRy/GwWIjhWdn4MNH4M7wUUBQ33ukapKRN4slJ7OJ+C2HmOe49jxjYLgdi
f2/iULlWZlt2njNn9ALlTsSeQ2NHboMZpfaD0vyYaCBz0ArHpU1Erv9pC5VXxxDfwp/kEHufACGy
uWvw8CTl94wMjjhTFQ6t2Q9D6MHT9HqxEpDcDF8fTYoJFPFUcJv/m/fYPNn1ox2wobV0TMejS38k
En8QEWf3YbhijFhmkG/2k/QH4V6NP53oeBhwdRAIvcW9CHRlMRECYclxEVjEc4yQNtyi5GPyS3Vf
vDQTPi7J7GfFJWGYClsMRvsTYXDCLegFnoV9/SoclzwffFYC/MRYjUQIBqQCKTUFYmS3H28dpPNi
68DRNlwQTYeAtQesBXOnsiCG0FgbERRdL4NzjO57wVcBPKB8skR2PwTBvX3bb7sabeiOcFs/EZWY
KO5xib2O+zB2ywV8yfhwBSe7Y72aGuMKad2k3iWGPmoqE/af09AjDX734b5wfL6h3pkzLx18bL2a
BKxMiyym95RRuYa6YDgisbslJem2XAyu8qeJXkwwmtcXs1lnQ9nAwbbwutHSY/uXjm1Wn+XWXeHO
yrtDhHI/YntP6xT+NSD4kb/m6dB12IwEg3cV8hLlc/RnBjjsBKsPWtcklBQwhymWllHy5D9tiPDa
PR1IM8rFpfpbTsuk7TKC+1U9yVy0K+O8tL8bu/Y4qBOtJ2Lw5ZQc3OkFDV3Ht+SawfiSgk7KWRlG
lEDw7oO1Ol4mrwHShe1fQy+EMfB8B4ATlKAqGw2L9kkBfxnBk+0Eeqg+x2zCdMTYJS+vvfMiMEu+
4URy4Lkee/Y6z/uBMSEWk0wC08YNUOlCqAXU2jCQ8iNcllXJVTikxUc7BOiEoaydCUFtn/NzJfKH
C0sZ1ijx9dV3fVN1n6owdAYhqx4htw3gOXM8C0nLkhPz/jfZ4PKvVyuDrMyVsGvkGsBKW1agnmT8
dh4cjxFe6dkliUiy50ro/OjD8BeFOJFzxxznt0x+bEA0KtZ4v7okbBCPMaMpOI51Pj0bYkpulLKt
CHrebJSRl5dh9twDao3VUiZ33dkKSPqRTr8+c+QHFTvNHz6X3FLR+/JoAEYI94cILYYcycFSbaMG
JtoDZjngoVDT2ox41o9yqT9ndQ7SAyAMFKm4akkOuBBQOy2NDMfky6vZxUXUv6TnPYo5ngIqfjlI
BBaYslYX7U5nCZroWVzVv1rUpgarFEPxwhhpHOJYq+P2bHofoGuvCQvUpQaHnnjAYn60LYtIkuos
O0QrdKaqts93YIxHFXShEX4tUTz9BTY4ZAO2KQK3HzElJKn6sq4LP9/wi0H6esian9kXBfAxhOnU
dbJKkqT+XClPJZqEwv+s2jx9n43wOou0q7aSnWNo3r8vrcQgSDAjh8tv4V+ahdFgapu2mTh/VGjy
zHCYcPlealnOFFyfB5sfPY4zkuwBk4QQr1/qPYN05LqBELe1qVadY7KjQ8lR3RySzaOmCb9IDmpA
Myr3q8lCes85CR/kS2KtVtEVgWzOhG0e93vrxEup2dQGSaHnPgHHj0RDUlySUZ5jtrM/kfX2kGGV
GI9sdEGJyWxHwGoxsXx4gXUG/oF7c/upoxZ0ap0oVIFtW/Jpu1yuLu5U7YQowXRc4e+jM07nPIpP
S8sSXTbfnDAdapYUWyVsHSg7dJUjbJN/YtSj9z5xiblFVO8QT++COQKpqzdpou5JLpEOPqQcNbJX
sys0NAseq0PEYLmZGwp1bEGYupYT95rb49ocfs0b6l3rFYwS7D4xRWh9l+ttswZtQpggWySDCvV1
bdZHTF+getfT3YBXdLnF873cCGtKeUYQBFFD6mRN8nR2KCDmpgZYhUwfBy+dVAcqhZedMQXTxKij
svyJyfiuxKUGgiWOSthrsdM3gSFOTiiZPeFl62kn/2oDjLKFfb9OaOLoeQ+y6SYLBQDdYWUPv5NL
p+n1bICX/8gQkGIEUNJ6HBku3NouKhVQK4Wbsr6lN+OuaZ8/y1b/FnHWk4Y8y75PWwTdjO5IvHS2
IAqgRrCaQ6LRQ0UE60n9phRIrI1pLCSzsRUOAgGiOOV1Jwa7Whq5yjkqEc+qQblmJIKNGbzABw8P
VMm/gsohzFR8fWY2GxOniFYY60G/uI8ad5Hd41C+QVKX1CTaV3vCf0xCu2vjCr7zRIEQaOxOLL68
qbOPXOyzYLAepBffHqlHkN4U2lQ6bRSyE9yS1NQbVRYcun9/O2+NR/+WVeiC1PEP0qEUKRUSkMWE
KIvdi32ilutlGTKsdCK6iyFtoAwi8CgZRetbCYf5hVwgnFSXRFPW01ZoWfUyYd7uGPah14n6JvGk
ewwjF0hcBc05A3P+Z97mi7zD+z6wqNY6ZLt5ULG57+tEd1NrOcVoPzAz7vHqjcKlhrtO92xurwIo
yi1Zq4ixBt7riRak34wbpT9fbc9bbRX+OWhwAzpq/XWwwj0omFv9Qf3IZBPa4NPrUFof82LxRscs
goEMdXBQtkG0mVh2tlFcaLVRWt+kainIT6r5+S9jK5Jrhy9UT6PMKIY/k9GyFQFD3D4DZF3BV7IZ
XKJbNbpTZxWYqlO6uJk6/FYCWCZ3MGk5YHyr+5BD4UGpJhuG9UO3K+kr0nE1q10gjEI8OTtSwjVo
mr19CC0xf0Ph+0UKSJkYxe6aPbdkfpJEGxCK4nJs5gpIhWhlVIx+oktyNE0qyAGEU/rpGXazfOjh
eLxp7Xzl2aIglFCd/6ZeLWZwV56GLlSUc4ux11t8rmxuKrbbaXkCKunQXnT5ySfwfe4y/hk3tb1v
QiSOsInhFHkncQ5FuCPDrPppKa186+p1Xap8fNXmdJYdQ2OhcT6XhLim8d2Wdt10vkVa2y2IG1+Y
goBy5/tSkwkao2thIE0OdSCjAyZ19mE0WrLacaKmHBD+hjWmnTPTR2e6PMYkpKIx7Nl8CQSOiGu2
9KM4gIkI0hkCzhE2sSmdycRQ7vEsDssM2Z+lXQVYZiaqYc9NoSQsxWdDHeNHlXtqbpIInXU4GCz5
NZM7Ojglp1tFC26gBZY/nTFAL8g39kIpW2GiRe5xYjsu6smEubABezWwQIFobLCg7kJV09O9a6qt
MgWCL+2+V0uKWeIzJlUqbkSoF01BAg1yEKqXvxGA+LOdvSFQjzo2qyTLFn6XzvW/KFKXxDDXtbLM
tIJKIlFI8v5j+2vkZD0Hup/bxj3y6LcOS3yeRJryfcixCp8Pnwsj9zYhpQOruQf1P463zvTgwA//
tiNalCWKuHAPwV028vzXlooQd42QptpdhJMZ9MB6Qx6K96wDl70Sw6jNm7nh85rtc4ZMzX6PnOXf
g/rgROJWe7Idimc7CZGmtIPvycl+Dc3szDuXLWRMAqVWV7ro7tXDfOt9LhjAqKM43mdYQ3/B1C5g
SEvXX5ai7LkFsSK/ZovLa3Ndk2vPSoLJZkAOCN6JwX2x7C8nMiGx3zc7wdTfxPOjrPDPTVpFaMm8
u9trCGj4bHQwZmETkRa5rhxXAHbr1NCLDcP8WM6irnUg8p9ijmiaZM6tdbU0ccZo9tn4MNvTXg2H
iDsWsB22U8LiOQsPe9DmoBm8YD0WCR+1DZXkPFXMRH8/zpucXjvaQU55QbJ+Gt02tl478YQNe72u
hppD837YGgLBVKeJAQ+wsyAtUQM/dlImc6fzUITZT7yPCWw/Q+Uhmtu1t+bt9cuxtpu0M6F/G11x
FnVcroMn+ae1PVkJRfPRWyV7v/Qg6Xrwvez/8IYcE6Zp0AQG0icdxZjBu383Gui+ztsr2EOHqTFe
s9N74AXFhKIJG8Jxo36QxheJ/LiHE3gKWRvrbeKaZRxp9RBh+5wUfGktDYcqxC5rkDSh2oVu3gFN
hTCS0Tpt+FbeJWMZuAPo4M4DNXxvuUV/Sg6ATELCvRHaPTVY9rlgYkPH3At8PArJgsQSXMii1Hgl
3VHTEhrlJrhmknrG6IIK4KmwaZDavVRTdACEzZwLdxPv9XjGIHA1gEKmYyVNxUeljVoG7XA+Kfdh
L8Q+WOR9JznvykEGopGJWARVzXiZOOKUCE2xKP3hRCS2mnbQ7C6z/3HUzX2KIV6oo1PzRZgV2RYB
pG+sa8Zl3ZXd49gLk++nwqgRsZd86cgXCcM/O+IT53NU9afMZ7Efe+33OBzJNcxzut4aH3ojEXIi
BIrkNQa0aJnFQFnGcVBQHq++czNmfz4iFv/g/TQB13gXzx3xvXRLaty20zZOrAKm2X3VLwBHCCBq
eMN7N1wz8VM8UP0UPv9pW7ZpDE9YSAyoERHdcWn8tVfrHO4H/iPhlEaFDUatEe9BqDEl6Mx4RK6i
vL2W4nL9iuL9uPtAyCN29W7QQq+ydWHpELTTA6jZARF2GJRcJxmAfL3XiS/vs8OSA1SCMChQwjHp
P7wqlCFLxoFszDGknVThkPpyiPJrcKusD2BKUqUv6P7XCqv+oJ3yoLJR677g6rcAgTtPw5qZmXVi
T2PG1U1qCO3/hhnpk8UCrbOiPILnsSVl6Bym5HuUuIGHKNX1x6sq2BxEX4sYwnOvbDmXntdqatSI
xG99UQIrbnRJet2pyP4LXvnPg/dmcqz1tyhxtFaXLimVh3XP9ZqSEDExjwXtiKjzk5XDQPGrbAx5
fH+YXcBynmih4VFekA1o4TbiqwfgFzYcGlC1BEV0f1pdPmr6al0zwUKGs3uJ0cmZdAfdizWebX5Q
q6ZVVttp71j8Jfdojgt3tsnrCnrwe//BxcUUmEMNhQU3dAPRg/c6rOPtCr9Upio1qJIP7cBw6WDQ
sxmxVgfTOxKpHsploMCtlkNl8cqJpfthbWbk2ryhIMlVkepRz/ROBeO3kU1ihDIjcnZhcNc0rXK6
hxk4Zub+J+dr+XpbFwPVeoZU7WbL+CZL73gPEbK0qpqdrBsZgE+zCURTgLL5IJI8c4bY4MSuD5d6
TkPknns5mpT52+44c9/lgPIadso2xbiaaJ6mZ5s3EiPh7JRzhKKzcP9hY2xRpKnIEyVq6HOvi0jY
UCQZ+f1g+mHuFsdPYeW+iZHhcYgbz5rAOnv46Wbu4+lYmKNKq0aGBTkoTtbmrftWvuM9pd5qqwgG
ETbsw1gqWTcENOgoWDeZNFjEAoEFt7bUlYWyGJVsVS2S+ymgvbnjiND7uVcn6SNva7lStwKrluJ2
rUY/Eg6ltyOZ/4UrW7dmmMH20/GFT5dKz8EoZk5nmXjFhIb1NnFfbX2X6AuYDVtgYLzirtnOAH1x
QbkvfzezQO1tzVAMGJMoO5YQ9S4jwf4yVxAUq1Oaimib29OUW5Q+QshzTyhfp2jOsE+Ugzwkfwd9
N7h+scXl8X5a28tiCizJNrvZ/xwYCn8A9u/jXevHPpm8I8F8q6mJzZo+Fu8Ptb7ZISO4pfLtB0Qx
dq5eH/MzWKH0Chx+9TqrTUwwTjboxIC96gym9BvAp8aWVTLWR3y37L90ncQDqiH/RSh/gO4Nutlx
Feq6sCt85DAts9lN+ZgQxUO83bizX5ZCoGrNJZOKowtLDDZRdlxptpaWLXHibBX8Vc9Vrk2L3Q2I
ZqzGnr6M+lZEK3VzrNcwiKu2rOylGGs88v7gkp7S8rYWQmJc5tOFJlEN6guW34HK2+24j02MY+Nz
V0iJHmgv3XpHpiVFBBhx0UzC0IWV7O0qn4KRtfHg9iq6dtQjdLar4wba9JihZ3L7sl1JPIOfxRm+
8rFJhgll0edxd4eak4k1qutme7T/tZLD0UG6ygX/dTWbsxEtqYZBk078K2XEzBSeAS7wl6wgOD3c
1IU0pXASkWfhnkM8BQDaqwcjAbUcF2kmgH8ZwwdM4h/KWc4LXah+dHJW7RJQf4SRmOIDLOYe3eLq
3Nho3G3lThvDnzb3DNcLvk9D6kiXiAZGKl5Y7g3v4zxSVcp1CAuwDkcxBFRx22wCQu9RNvvyAS0t
EaEK7Ace7DiI4MX5YsQOY4tA36HKmuNgzMrNlOBx8wvlwUWnt3ublOjfuddfoditCMpgBDPPve48
g230eayjg3QxyBtF9Pc62P0Q3CJXyUAGrzvm7yBLIW6/DTQ5EIWcswtmZf7jfGoAm/p6eZbViGPp
jI2fXFQQXWqJzgpf1N1OTuIaaHWxNXmvFTZuvFvsoSRFAxU14384Yx9lrpOlDVzrgZxkQNXqgMyH
XGzUi3hTY0/i4FmXgLo/E8+iRzfEiYdAW978J5IiI388aPU4xkVEGLBraWu+dIXese0K3/FXDF6C
dCN9UoHD+QqCYDWSphsspLxaAG9fwvyhsXHgVtfdnAinqJfPWXkn6T4JJahklJ52NVkEODmPuKKo
MKSW5QjY5fvtLvk/2vyhTO8Fy0gqZw3wbVLdVCRwUQC59EzPTH0AH6m8lYNMsLVFtkSPl9fGJBqf
98XcLd0B+rcOvLHVUmlu58q3rSTadlJlUfC9/KITQy7NttQbPcfvBnnFkutX0Sh/43Crd/w4x8h0
DghIZzr/4ZdHIrwQaqcA2Bgp52+ZVwoxUAyZsZDCykJoLyE8qwJUKewFeWlhPA4eVG5KUQob/fb5
KXTkSnpbUdbJNmUncvx5NUkGTdB+KbTKVhgmHIdrZ04vl16RVuv1jOtvrAjlN8ngPDTkoMF4V/gx
hYay+LrvNInVaCADn6OLy3iHAbAdlnmUQVitFD6FQjLmEkK5iZ9DTPFNnjVzrQHacwYiRN8S8/7t
3vcNxRsm9Qk0cS7S+j5vnr5pnE92jCM+O4Qt7tzVQnYb0Wfhr6REOUj4UKH0TbL6A6qV1+MsSwJf
DgEdGrHrD1rWfsway/h3YQIio6k9O/0KdphLqBmGJbiQCZ59d9OC78QPFYE0hIyDvRJJKsmOEQb4
tY2J5jc8AuVwOZNDjMN/9jWx60EcRppURyaDTj4nUGdzXftRGdpOPwxzCDIe1DHpwZRjD/m/eGpx
nrZxFZo8zAuizKoOye5x2lL23CnCp97tvj1vyDhUtajz0ze9ngy/lQYT8Lvsm+f6QtLK2j56b4jK
0XD9EoGnZbWfC02mIy3OQ8k1KjC1c5/qHD6q4LEscSYxujyvesg0LWIXje0fpUGVZXZA4gITb6i3
SQrSmuTDLLEtKjAp6b9FMcDoavdLG86fOIluCx0+6D3GuTn/v+8Bi98ry9FlQ0PpDn/fj/xvyUAQ
6nwpAYYHUy9eZ9Z3T/QHuze58Np7RlhH3Hu1+Ok7YkZb9H93oPip8DZnQZMmZwMdVER/ZdPE/oi9
EFTariFkvXsoW0s+oZXWvVx8s304g6xTGjVfxmEWyCyvcZbNVhyI0J2ay1v3qiczFDWfG7yL+rtW
BEV0Q/G/qwWE7OGxJIVmr/Zc9ngQbuEXDV9flj8l4To4YLihWwMVvfDntx5gxGaqlJbWsN+tt6qi
4mY1AdJQYttd+aTFgzgISrugzw7m2Wk1Hbw+sjy9j5oVMMcPBNV7QWbndDiBwQZruOP5EBB0Cons
YgKmMPEdb94hNyhgt3xFKUK4ifsZ+FZow42wnUpPxNvsq9ttMX08p2SiliUqI0nmMUPSMHD3/b6o
s8Xzj+uup0GuW9kec0tg8euM/A7LIBkbq4MmD1Zp013Xy7557Btlc/PhGc7V1XXnCammCrlXCyvR
4Z8NoAl5TuhLrDcZcPM9/LzAeY1KWx7ec/R4jAQDSD6bQpAWNuLooP8gAdTw6dULiWgDVUw+ATzj
e5jPl5vhQCtZwLw9CkMG5FTa27RzOnffSpy1AE+2U8pebnlMCVPe+RpKMg6p1vRj/W5rBY+iCPE5
SXIKHg/k1K1tvoWdcyRGdpd5YWpVROwRlMddlMf6DA5syG1beRsg5hyl1RFlQNAp0vrYaYs0u4Vl
+i1yEyNgURY4WW1j7PCywsNmvJEkI8Amo6LFN2jzFyEoKj1tOYm5flNLn+JZy75ILeyJ0dD1PjqX
+Hp0YCFhKaReiZfNnkLXnsOzCu1mRBc8aiZ3eZ3WtajX2mJLYbZjbXLbeDM8RMSjyODq9SJpQbJj
NS9mnouOgCyhS5YZPBSFpo3q1v9tthwNrL9CQZWXd8IUr2YTDK0QExc80U1EfT44l/pa+7W3bxJA
FAAJdSklw4NCZ8kTpw0ySM3HHIhyTNS9e61fGghifT2CG3E5Qz/w0nj0rYdR2XDpHZzF/2pCasOg
K86s+dY09ebrn6av92HXh2kT11U1TRWDbhGzfPAstxnA+fEU5u7suTXuLo/zOpDQGf6kXAc+ACej
ibTF+nDcpqLZpb062uSBNzg897ionDE6EAvBiqVkujVCCeWfTw98hgsin0DS1UfJTI710Tki7hxf
k4r1f/Oo9/bjA1VbRg7hMWLxhVyfhX12LryKxbmlkUk0BSxxB3hqOYZycNXtrLOzg0RvsF0ksYmV
WBiFDGDZirXf5DZzYc+iKerum78zlfoSpK2OGE7Jc1qF8mXny3+wJjmp009tXvt6SNKSgicPTHN2
a/+o3+gqWBX9g+Yq9QYy+Mzr/72I5+8jEpm/QXtf2yrYb/pUd6CbPPjqDFgimbyhVTZxxwBh4ozH
SqoZ5KZqLClNJm859PcciFUwwLK8EJ6mTDDJUKoRANOMR1ktkCnoMxMjkptxKsGzcXQ+PtykSYzc
6qfDgPP7AiCX8+hXOs4kCQEpWE2MbvsBZkuc6ua5HvfzxMTX6YguC8tmy83DRF9SHqfa7imlTZd0
7DB42g7vVKAwriabTvvVCjI8qxay/PtpG7MudhvxEYtx3TIIe0nVWLAuYSXdoAL3Fd2SwCmIAilB
InWZxaNC1uoCUPpCJJwZgCfVLQHbiIjs0skLUX7mWhf7IqmwprYFeGTVm6I8zot0ghC48Swc61Tz
VL7AAXVKRRItSNJIz2yh9sVW1PVfvXiOvYpQ79VUB9ai4txKz4icN4cngxIDfjlhNQzg3Lj2oWUW
j3fBPaUy/BYGFki1oqiAh/hJf6EhE13qJ5hfTE7vButOj2MKamDqzSnJmCxNADCW2W8lYGVfSNfF
cycZc3Gv7P7oYkiPraWFITrS+N+jjx/BvV20270ddJISAXsp1yv/X5hRHRrvCKt3SuCpmAp3lWdv
2enqkHvv2aO0UH3RWhC67AllTPfKimI1TJM/22AKELynokWbv/xu3NB/iJlm8jdcSnbNUkZGNokV
S+X5bhPhxleBPUpekt90qaiDPnuSr6ohEzYBtdbFcnAtFmyx0SdLeuYCD5Ke4Xq6OvTK/FSw4YPR
+gXEDk7DmVUg2oX+ceU9Ry5j2rCBhflG6IMj56BCV9UZ3HnrS7BapArI4ajX4vIYeQTl63lq2xZj
bJsVG5w9qDmepnRzCZb5Jznl8dYHRFbIUW3odqaMBBv7aTNYnkmfTBQ9v/VNtOHXDOQLk2WR80oL
F+aVxdGMxJzTlRCTZSVF0uk1uwD//rJ5xAX4XZKaSi9kT9A4YR9eseE6Gd0dnxY6PgNk56lBofQU
7fvxAMrshI09PE0ugpPT152LxdXtJjLshIlexqf7CpMj65UFjq55I7EkaAMSzBD5s67ukQ9R+ZRM
fo8IQy/vjkvwbtIemwYUgPlfr+cVaDJlnuTIxAmNNi+IqWuUKs4R0bpddbP7Bas5R77ku4wGgnU/
SaQO9Q4dz4dWsJInwSK3Ddt9SP96PQgCHbXbPNED4wJztAg/VbVh9RGswa/HwuccPwIHo2gg8WOK
b06EpYwkFAaAyquJOm19C40q5XkZBwMcTYvmhT29ybK0FCiQ1z78qTH6jRt9d6bNFPqhkW6zNXzm
k1/WufBIRN8ve+Cuu2Wwiq53oO+JB6uHI3UJBKN19zvzkTtlFUUS7cPj0LdQrl89U+OK/+S5Etuu
mjTQdd86TF1DKqmyJz/Cln2R0QeUV/zWDj0aAYFXk7USLglgCKu4/H0NRvyrvWkaBzBbO09yCPkx
ls1RAHW7fhH9arptrNXWYUGOv+abtFC9Y0LAOnhpv5oCL7aSH8ZlSVXyHrn6zvs467P0QMg3MWfh
6EO3VKO0cUXbtvqAHQNvm+yPrikgMJJpObTGd/oQsPvg4FEYAZCACWtLgYyJCagWqjYcTehEbD1e
a8icwbRJzH3DRrQR7JFeEAx4N69ZsVWeqahOU9kSOM4Th1zqEgY1FaVqWgrhXdFTfF7tE0uwz6+O
2ZTNxPl56eiccZSh6ihqAVtkwcg7A5qfpuIF9qpTaq1u2YYJIKQPl/+CoQTlN0XK4UmsrkvJWM65
m6RTQTW2YDhwdqoLtMQF5mK+FZwzzp4CrFk6g4gW67RhvxggdDWtuyec1VNO7ubisWCxY/l5/dyc
WGnDL5TwCxykYynEYwerIhucbgNeFQtpiHnxqsm7u9iY2nb6OFZBTeyYxW+PfzXR7ijkERrs+5At
lJQH1qryeIL6SzQBSJQXwGYE+cvyabpSLPzbCGbjpVz8KM3r9dzJ88FtoucJfClL7ns2KHjC6AYn
NDsf0S63lMbvHqBe1n58eCybe+GV9BAU61s0zww7QnWbu/uNPF7P+RC/6AY6aR+Pz9FkGk6Ncr8b
jXYXNKbvBYo/UMuCWP4EyCQHzq7v4IvcbptjF87aUogvSfUUQXqZ6guov6Yhd07cyFJzsE+v582C
+eIMWmO3tYm7nnHLz7x6vDA+OydrKWE4XGruW3RASTdd/dX/knYsgqPGCbVoVl9NiC0fuv0Mc4IY
q9aOorA4l8jrO2me3yt5t4HTRxZwSybuLAgp1DNmcJj8AhhO4S0lEmP3xWJGRFi4KPc8bjJi3JL1
qBmEvMJ4wKcggG28Je124v81UB+k6HM3pdV3b8T5gIYR5RrnxzYkXD/brS2e6eqJFf2o2aMURhaI
WmkBBNlPKEK56MyM5kPdPomo8zupgviQR435+A/cNEdRlN1Elv+42+BvYJxfqNTugBOiW32058k8
9bNoO/onsQlvAACqrJZioXrAnWnwxFB9DFka6GGdruvfgJdGdvvUI2CdSnYggDYRUUMMGpentA+/
kCLOi34xdAJxK5AqNKJOM2oNQPpxKhy3QI/vu8PcHCqE6dUU5etQCdToLizA/JKQ0Nd0BVCKJlGg
Dqf0wfu1fwZTbFU04MAiKPHpJL8KxLCvzk7Ajv0l3cskQVD3kxdoc9lmwVEW74or7F/MQd2Mp7q6
8RKQ2Zy2tvKb20cfQ9EM+4u5Cr/OicCMb5PB7suK7lwvrG4cc5kptr7mgJhX3kd7ec0mI6aoXE5E
iKM7KcAvHZHkvwS38LglYMY01le5q8k8/COyfor1NCDWG90j1j/Z2FqT9Ne9oJSWCkOSFJbg0+Wx
eI3nG7za1wqaYDXXdKJW3rB/6HKHM9RYaWJMofTO+3KOpd2tg8UNawc1h3z7xDcSa/Fkqw4f7rDz
P7iae8QuC5lMmn1p9OXzD23pBxH8K7QSpE4ih5hDUm/ecjAWiFPD8WOf/TiPvf9Y8zAaJpDZ1EVk
DY5fEHTi43OFTH+WkutfrAj1vs/ABIaylyc/ifF055iBZ82yfxrEx41jR2iFKK42Cp1C1C5Flco7
55Qqme6eGf5XZZIm+nU9VYD0gSMdO13WUDSvdG54K6ejEgCPbvap8SplUtvZW2ipq0TUsjlbOxqJ
J3ZmhnuKw6CwbZox7j1Z2fiSPxJbVViRYidCaRCJn84iQkaiuw+YnHzPKGZyjdPR0op9zZU8PHxE
nl2qyaCeXkvSiOAhZd82yboMMkKaw3OwkDGnpKf1a3omtRGx1B3EMtRBXljuZtj9stwJ3nNKNFN1
lOiyXiWpCf4xPPfqpmWp8XINCMpA8xO0k1Y0ve2/qeb6MjKvAifY7dP6mpl3Nqiy3z4kM6/ux2TR
iCV8Z9j9sbARSangwZHAJJfmS7QojffqK6M/50TiXGLY61zaB7eOcrrKiX3njwpYzqITOlP0YAxb
j4aw8KFSJgHBYId7ygJzJhBwWLbx8UbXbtObfkUWWCbgL3+AhKe5/s0vxz8K7M2jTauw7Nf2o22K
JRifZreadTlwOjuKwvODb3CL7N+hYjqjL+ryPBENDJtgZUKC+jaIpgMmfKVbQkjOrL35jb92pQgK
cvtfKlodnDSreewG0DVQ6318xOF5N6p2KTNJxCD7Mp175ElahweD5h1TRsOVR+OfhnWLztiTZbH1
OW2clzvtVbo00mKooEu7XYIl6oSjiX+2R1RoXET997YIpiAuZ596InKzj//KynsG0IRdkpwju+PW
3jJTIHwCfm+Kp7hshKTc33ZGYYxABmjXf3FrTqyttF8b90lbUd5eRJAQCKgFnm2CRslVADKykU0Y
RN5SCfcqTZ5/KSBSeknENd0QUSpBLXvHpMh7dNJxxPn8VlAL81BHnhngP4w2k5PUHZ9yYWabOnQ4
gdQzvwGDDBUEF3ZGAB6kQuWE35xtFgV/ExEHy/RS7376qNY+TXL6Lz5Tjqsji4KeFy5STcUzqpzM
aZFT7DHKlM2ExFILeMchoVCCfradkj0w1xiq/HJPMQIlxDES20suGW6z/y0Lh6LJHVrNpX1F+m8a
DOUcKYtcQelNR66f9C/2epBxMouA/k0Wxd6N3B30TWdvCXMO6v0lwzOjgY6/Ekuif7xnJJabxicJ
v1MkAXH/YehxxujUiF3Fmp0vw/qWqyIiFuc7TXqc9o0urYXYPNI41JeBYN8tP9S7lfISDaf/PMrm
7NqFKZ0kz91KMyAtojMuFV968ONeQ+qi78L/6/Yz4I+dALrqnuA+EkWuKEq8X8/40EXBC/WJt+et
Kwh8JxwY1ZmLUh6dBOTMzhgiZDxjsTXXMeCyCrLa0q3H1rFzpPpgIZJaU/laiyHv8anV5pOiU2mA
vj/hrXhqs0qt7qOXA0svewA2DZgqPkgWLJWPEur7cACR9uRWKk4SveyCjcdYLWMLFJuehWUX+jju
LOKIsQ/M91AiLen9+LpQIhoOgvn/CWuxrQZffBLxrmkWs/WPAMtrcQ8rWINrPm75MaUnTcWg108K
rOUrCuFlVO4xbhz5grwUVfLrI190hX3ol/SzPuUcWvTNQx/CZXs/zxLp542VtUGZCDyGmBneYHLc
Xvpm+31eGvTYXEV3PgKaMM9++nmT9ANuM1iDK/6gEh5qqF0CgcZD5fPH5TxKCxsb22I6s9e/kRVk
pCzi1v7dRSK9CpuHKBCm4FAk8mBklDRHi2T141VW6siYEDsf2Acuul7WsfsMzy2QVSIrtvfUrO8l
yoNyTmg/HX/itcT1DPXkuv7Lp1rmGGttVBxiQj74dLaTknrSB3cRgCFFcdcL2sZoVYIVtTDF0qPq
XRqxLCTb/Q3THkPdCHc8fajB37FOEgzbFUSEYYIJCHm0OGyIOnfBFdOt5AtcYmWPRDAj643+H0jy
efsuM4VqgJZ7m+KPwtsmP81TfmGZHnqXykv7r7ZJv/c0tjc/gHqVLEIhyyMy3gHDpc1n+BVh77BU
x/RlKxyn9ZNH0yCzhc9GXC6KzbWa7M6CzGXDV8YtFk6p7fBqDtM3297Zn4q0XG/eI6M9yqHKH03B
8i9ykf802njdQa2pOG2gD95VRCPpm8dGEuAyse/FfkJN2NWus9FcNfd5OsGC4PrLukSgfqd3bsKC
CLbWEM7U+mRtwqhB2q5789alaHUzZmHcge+gR5qw0AOpMUfEOlRBCjJEMGHamvqxH5XtCrYdwFL6
nXg+9qeN+Q6AaN9KXrluOaepsi+OQDl3SgxNBcye4wiQEKfnySTsJasshTQSeKAIoRmORiXAZbDX
SU+oeVbVUrHbBhrQHSyQlJP579bcKdwRtGbVhpR3Nia8nPZdXE5mt1M59upVWt3qWjMWguq+sSvi
anWfQ+13MFkbhDVcfYWyil3gQ2V2H5ImSVI9Kk8QIZxc/7rWkA6tOjEA/0CfB5lEKkjp4vgl0aA5
jzh1xz62D3mvoGGRD2ijg5y4I3eNQ5GiEmZdDjJFjjYUMPWToYWRCHXiyBDMpl0m/vdyeOxFnb8w
09lHfvwtfK7/HHlIsjyTRMd102IfIrRzdkOuE7NqNAt3CoGVnuuRfhh4UIyE1lexu6feprfJ88kB
1EBfnsxdGNBQkAjeKrl6003E37WSbbUWvfbZtLPdY4yCfn7mOzcDIiZDGGpeAi1P9Ces2YZkME2a
jeM6aeobuetpgjt+huHUg3HseWlQ4DctwhKbb+NNfAcA+t6Fv+2E2PPGl/75E1K9sfvEIqIILSr2
clPXwS1nmHjhNLdFyT5OisjACBnXuAmXRWnrmQ7UQj5/pYSZgMt1pwzwaEeD9vcvjgGPnSdUBynH
EnR9HNyi+oLXkAiwpTySMpKlApU0ZAwglpMD4ZuuHJNdd1sFwwMyDIhwdgZkyZ5SZS9WWQuUQXJb
7a7kZGgdEzrnSiHsVB1e1IidY6oDPUtTHjqxzbC3j5oi74DrsadSI6VewbNTJwGZFVmeNkJK+gEb
eUS9aEkFTDZGF0FuthYWN/vQ9AHtQvIhXEH3A3PisFgNVvnW45RHppQ0eLCOxNMEJN145RNv8vZS
W4Lazn0EWHCZJ//zjISR/f6iymxTB5rjpRGq7xgBZv83eJlNMMJLDvZmB95DP7Q3px+ZumS02elE
mJ+8C/JvWfN++n9+dAsoQSBbhf7ob5caE0qCr2gXkDL7bzAfKVa14M8kixNeMoYcfn2PNw4rbwyc
WZbPNXibNKtYz4NIIpHnIuBZsIx3GygrjHqfPHcAikYKmRM0OzmJiSAVhpAg+MdfJBhQ0+QhJuNg
qQUVgZlzkxnKJHmXt8STJXDbaOvWu2McZ11sU9Wxry1nOalP7DLg4/0B2Ekx2aZTPr/DQRZ/eaRr
TMMKKkZKd8+keXTl8khIgmGyivpXsi9ayXuJSRijpdzgUVuYzwMOLVgvyiUmJzN/AQhjiwH76hrg
Y04bo4oZwsNWXG9z6bhGVoCu5B21oUNjc1Ur/Vp2STSozkvoYua8ZgYHmfvuIt5gu9dMe6alMscG
E5+fHJVur7yu4CTUGV8ATssHBaD2dwjWMqtwncZ7wlw9vS5JTAJBqbOJyboq6YOEscfAOdx45zAp
r2+7lLQ5iX3UDDXXAIFiF58gfsV+kJbVmtlHlSjFDuhQhq46sKXmSvS9Mth+lKXYlwkxvs3Aer4g
yso6PR7U47vdpr9RzwBr9//+5HAjuNciX3vuaGt5+mh/tIFm926aE23QSW5zoA9+XkUIawzSfUwN
BuTxChuCbBoTzzwJsAKDYPwF0FMcT8YtUv40effa1lXQLkcrrXaaElifqi23lk7c5B2KYigSsrx8
1kjG5JuHfXDRNnZgDcc9C9WW9crErb1ZTxT5F9VRavQ4ISg9H5eCjFLDWuxkb1fxN8ES+NfcgT8f
GicUtHJHRKN2YZx9qamS5vtsj2CGor2bEhYx81JX8ga17mmRniWtBjkzxXw2fYbghmNWsY+USsf3
OWXIoaaIRU/XARAcqq441h9EFz2457nwXrkEfaRhg+KU7rucy3nFNokHBBgBi6lr3MLQsUJ+tyPt
rGQwWNNmbHzDTkHq6O9qUK3stvf5qyn1wuQ17yhN4v9efJ+TVwoTJB3bB0kRr27aKRixTZJ5Sb7x
fAOds+kqgcAzy0ZOXwToUNY4awhcJD77gw9YBnKFdSY0c86WqlAzfbpLwWe8yVhZly8Rxis3l/iw
+snacvFFrkm6982ZZrP/aIKmOerqum/az24GkZKYgnntkFoW7SVxYXv3/+2V93PAA5C9pum8qE5S
pY/tYppaHgfRiN7vApmo2g2YNdi9f3MEx51HrO0pdc2wyUK5Lg/tJ0zG4vCCO2JG/AVUm85I8eE0
EJY4HJDFnUcHBsKvB9RxG270oKbqYMpD7C1LQ+O8Pxw6Q9/M2xq2hnCs5cEWJe+PJbzSrDtOFF8m
3828KnvBUsXuiZxon0MaQZZe0m34QbHHg66cs0lx3KA2XNw0INi94oDCqEk4M5kAV56Ej2poCOqM
quEUJCJqlsJc7u0e9wI7oItcPTvzJC6S02hLRsV8xYcENw3yRX8ypN2VLCeQ0cCLGK/Pxv0gvCtQ
FQL5R9J00pqBiyPmIE5X3G1JPniHjshrIpkm3CQ3Dw5PPDnjbB4dnD+r6fBiYQsw2OE1FZZ1kPZh
xyKtT+y9i79Sx3y5YJ4M9/4Dmnrem7muYRgF2sMc3fhDBDSAH8KrAE1Tn4jBW2iTJF6V3Ml+6FK1
iKjiHCsxr6nyg7Lw25PUG54n+Y1o8axVMN6BGVL+s6HsA5PomuJdBRsiOb0BFqx+20qUG/zdKnll
jfNpGlXWKQ0a3hoJEiCtG0K50R0LQe2ku8Beb6/1PEUg1PhGy+1d2VDm6q4Kiwe5/1jc7ByCWmgv
aCmNwVWjF1u/RcvZtdpQd6vWMJmjXlecMuHFH7Dnmj2rC8OUR5/PDRjFLvij3pZStrwkN6CQ9HY6
AHVyKCrsheIRn+zfbbw9cESgiMT9o0bnpnFJ+UFXYVT0b5gO25DbEnyt/dglSIHgXQkUinuoBreC
6F7/fUmY4k/z2M/WSxuqKLA7Mcc1/Lac8gyErX1Lz3iGItCD5oZFxkA+Q1ftCW3cKigJaHLHzfVG
s4D8w5AwyguaJJrU631bA5HG7zgEckMf8kv6ORh/fwLT5TwxvloPf6oWSRosTavlnP5KTN+udLFZ
21yITwUuBYf042KjOPCON15U+BiAzTnuB5/edxPE4Q6l0ZW60TEJ1r91pIus6iyPYuLEVaaCyDCn
vCWlZCFTKVHcz61p8jShOYRmKe2ZrJfSQgEsMB8oeIgnucjj0rL4Xg2CqoGamxPj21JWKc/NAxrn
FNTI0WYMTa+pdn462RAdpNfWtEmMha7DJtszOiDOb0D35ziIx+j1B+6eyuV/QJ0PpQahoBR8Qgv/
Wwr2sAZfsnaMG8hJufyZeZNjwIItgEGrJB0PqhrOHgf9TlgsIQCaYBG4DGsw22LFLjgD6N44Cllx
OwX3CK4T4rKXyNKI04bFpBJ9631xiO0HyPJpQJv5g4eAKjR8BgmxaoTwF364uGIyLzlzx7FOSvLO
HU1gLrW8Qd4ShlcPoeLT2q9UEdjjbc0ads+cjlx1EjtBf9AI5DsO5zpE2Sd59oncIFRgEboYg6Wy
lRTRJOG603GzZNwrpVJarmz+nly1sK21n7wxg10magFbBVkXwDkH1WwNaDxOa2YEKRnP2yX9xgPH
0gyPgz3L4zm/bMU+M30N0JXbLGsoGM9dSS0wORRRE+2WruC4mCq1Ch4GxyBotVAU5HX+hYPWL4oC
tIXtgAY1MIWft6jkpMW92kCiNnBGRdmT4uDUBwUBG90fOB4fjW9PZIL7MCsxLWkOlZVxVRYEal/V
S2Z4mfigObkowwz3VseVShck9jnJ5MLMoCG0f0DWguPJEIWVyuFpunWIp0kOdGQYHPf4fQui9Pep
oWLrLvS7jAVDSG+mNc4h+ZKq/ubkdaIcE4jI2B7ssXrbc1bY+ZtCgsMCZhzfpf+TZA044ZatqAWo
dQYhmzFVGKyfc6WKfjsaOfT1gGu+LDIKOxop71OCUHTznSfGXFoCBPuPz097h8X9RxyzO+o9BnXS
2Bi7lgy9r5fgEXU7+DAr5bm1Dk9sOfBnJY1kgAsHuo/rx9UiSToA84lhlBSuU6+b2IhsGxpYa96H
/LveSTVO5riJ+wh/iFpfDZIFRSFzDLQUILX3JARnPB2tbZDu+e41JBxVBuiNN4GL1AnJgZ6ECKCs
YLeug0iqC+3+QlMAWdg5pOUBznJfI+WhS+zcMV7Rj2k1I7kjeqonXryOrwVruX5bp7bUpv30L6Hx
JtP8xo/hS2fv0Pi6bh75QYndvpIZx0LRMdeQ6UdHBOyKtHWmgbxdjFt42L4Ldc7kQDBR4Gb5Z9Id
S7YRKI6DS2NmUttpJwzbkB7P/L1B44fcR1VKFKk2R0vcFuKTCEBv463ENfJZQKucQOJHj4Fv8MK5
nOnsMONGADAi4ATd4fGsGE67fxhE5PVAzoCYKtNwHSf82UW3UFna1xPJUWDoLKkG1esc9ZL00v0/
yTN1HhdOMdd+qhet6KbcyCQxWZnjOsEhgGUnawC/mMQ3aTDaISM+skMSHkKcu92jjFUq0GpWnWYV
d6iYLTLL9tXR9T/8Swg25iyzRtn+qN4l5NzJPgHJp8rBiofvPJwP2OfAlKMkLxIhwBlgJG8Olxv7
XqmiVUXPb7AmWsnVoE4U+R9bDort42bqyP4LF8h/SPb9Xl7Ng397+7soZGSH9uasVdWEr0i3a5mk
mWCTyKEOwtt24rTDC5jA5EcvQ7x6uVRGWPqRllCsojwcEjAS9gQ2HPD4jSYZbdgUsP+Zs3vHXCRY
3Hdh3wLi8dYmyA2+b4+/gv0ChIjNHIqUYiPkjaOgLKs1DlsEl8GQS4diu4I3rdaKtYdJi1hwkiDX
VbDJdyO/R+r9Cec8dhfRuwduxMXyVa7I7PT7G/z2lu66NuyyTHP4EEqXdmv5ubS/6I2u0FV67Jr/
bPNMxlbYcV70R4Yp+O1cAoKC0JPXn6LBXVxti5VVlWQoVQphzyPyZRvGq9BkpUwZsQOUP3wSy6Zs
JayNkhSotXlmJi0/a0VIiNFZzidzbP25u6KoQzm81fVAZBHOwivMqNE9HJWj420iJ/WEjXD+lc2K
rVc2vTxuYz6bj0T6fstcWu6r/A13w2nsNZuhyYjeUJlTKAhgd56WPbZhmDMyQZAbwHXa5AKSpnn5
GKyzuT2afGgnvpbyHUYpIjcFu38RpUmto4bRmBKB83m3IdoiWN1XxMD/Yx17k8ULUfU8JElbwU9x
5bnDFRMLCecSJmtlPVUheinmD+XayCX/BT7dFOqovMua3xpmy5/bwjhyUJ7kQGf1yi9ZbaMZnOpu
Vnpt9TdDBbZ1LtXIokqmpWg0LFBOfZah+KAfZQaL1cQZssg3qRJDRRNy8gapUoUfM8wTGgkFci66
rtkC4YDgNg88BctphAjqNmZ4cUH8tzG2MGyFhqpvOhmrkl/fb6OH/7Ak4jqpIttRaUthyJQzEmQM
xfsWvMoBO5VB0hO1zdf0+h5u3CE0b4G3M2p5xGIQQXvb3UoF1hQihWcPWqCbQDuoQGFcUTJsMm9S
s31G3yPe+anx/eb34rKEl/u9MdwlyVlfm6TdnYldfzhv9EU/e6ghlzSPmJ7xxUyH+f6kcsVKS0Ox
w8gaMptcPkt89TnUD7v3BeZNfTZ1KwR/S/u25T9LK7/5dYTAi9py1n4s967IkX5OcKCJPZdHnLy3
/2GHUxXUgACVv4cXuvcjt2HoDGtVN/KIoLY6UD+4U0m8nMs4li1jjUZjj2wJWCLHCfhsdKvtkKAy
4O21sgY+q/XYPyw9mEstBwB4kfXlrohndCWMoP1L/f17MemUde11iTgwyXzbtLgLoh6Ng6jLVnM2
IzTDIqFXIeGRl1oJTXlRT41z3A/uHmLcDnNsiyVo0A2NwpnoWvwLAF3L+M04rjGuntHc4/6ZWviq
bfgg5NVNOP4ytLEqcsc4kun8kpL0MZ0pxIVWk1ly6zuhGxizG2KS1kw9KTw3T2djE+bnn8FrA3pH
DPeCBihk9FAKOuBoV2QH3fYU+f2da3Bwh0h9Imp47i9mZagPPgsPRRDCPQr83cfoeln4Cqfn9DXv
WQlW6bd8Mf0kqi/YfvEzUH81/Lk098FrdMlCrrIjNsHM5pPnKy+MsmVzppoXadUUt5+iI/ZCt+Aj
DIbAX7Uls7U/X8bkX34ZekjDhNj9Bch84dFw3dqAqNqmGiJfpfhzx3n2cZNFrCY2RP6jfG1cRX6t
+JUnvfbbc905XokAuH35/N9XDXxgb77i8U+Lu33ga/pZCtR6WFTaDNLDYTiqMUksvaYuhW+Sin7h
wd2QJlgo6CMqqTXBtKRe1+Y6nWYR8IMaFpAKZsWpKMHx1gxHIuZsWvCtbBXhF9oKVusmdjAtgzXP
v6Fhw4kY1wezAlqn8HONf4B6cYYza2ikVOpj11o2eM0DykJ9nqePuzWITBr0tGPjS5NAI+LOU8lH
nO6g1TpKMR7JmC1Rq/+Eo1FZTw7CoL3tjy9aFLyajgwdjkjFd3BhEKhIAPJbAjYuZwojpehrh5wY
+FAfmrN2m2vA6aOpkR5ltR8Fpd8q8fjgtna90iKVf6iIAxt9reaQX4DvXmmCGho+YapeBCYGaA/z
pY36QEo4sf8n73AuWf675s+Br2MVeNFcAifAE6mIP+IuqgBLRzPePOGc0pFeiM9rc5VPX1H1+aKq
scTW2FCK1/H+4wCkbJchGNw/TUoJ/oMtUaSa1xB3aUsKu6fsizCn5phJykLHSHP4Us17IKC6/QKP
LV9Dsb5oOW07XnBWBwW0QTqKhmhFMHRE96o7+PGYuO8jVEkpAux3yBw44+b6pfMaiB1qVZXSWYUu
enhwKQzOMI4D2U+6chXiYTuTbqmOFjDk3KuWhDzDEwK7pQUAAUMoc9sQEf0h8qPGvDMbI5zmWYES
IkzVC80wXbOhQ/f65xerntR4HS8Rj62nN15i9QW7HHN/Y6flJLkgFS1mFtJjrLwCio6Tj1ZX0Kfn
xvpjt6izvCIh+5X8pg7ZmTtxVmg4nApKOxedlTHZq9IPNYT2lkgX7bKnuNRDg2nUY+Hnpl7oYRCa
o5qE+f+VzT/mTsGucT6vvCf+PhsFeTajfhVcEAmj9uaOBPWNGy32lHW7p5mJQykbHHvcm4Uov0un
rWsjImZePt8wcfHUC8FMUXpt5EvSqQkUtQ52QzVE8GVmb61AaPDVqH/ZH3dwWxJVpHC8JCjlGjUl
Q/hh/N4A1NcsInYb2qw6NFgXUDkXqdLrtHiTuWfLP3fLyqRZJbCiykYvV2Ag7b8VUvkydcrrVTXA
GOHWwBNIdqqNszSm0YHsQBde8fBBdKMiqRXq9x2U/z/2jIm/taXc+yMM8jzNLAim00nav7YXtRIH
XtNmZkRlko1PFdEafaDNfXAQ6jTjia1buCAGRi0Nd+oOhSYdgCBlGQQuMkUh6hu17akveBi4MJOn
eynxvRZSZayH5DweoeNuUIHsdeTLKR7MhCqapvzJMAcVqaOzgao6+Twqb2N1Ef/b5ETR9OH3fHTX
6yhdl2yk4stVgeNcVgIJrRFKmesfwCosedRCKQNzRQIBAV8KqKmxbQLAHx82tjriMvBM3dbU/kCg
zQ+AhIFgMFv9ME+ATmhyxalkYxBzZvPpeWogInTgeOKfRenqVy1/7EICNj9MDhn1Sf1Q6ew8jHY6
+gNh632x8Q+2Uh6+ywl7RjpjPu2WJGlN31yDjK/hgbx1LJIv8QKRjdwlGxTSeBRhM4luvgubvUAz
0WUnk5O5GmRcIg0r4QVothvpYy9+18gObgKRcArYnkqI4OwTTDH8CGVl15A03DFzNaqHLdNGyb+b
2tBbz1mvl9248RXAaMfOFilXu0213dfUV9Scrlf6r5JNadO7r6RUNW7aeGO37DcEoltzHLtHVYm1
EVD1jyR9HuJhBviUUj7jB0ULBxd1A0rqiQGo4C6LNDc7WaD7iCzuF6y06JVlqHb3slpj47A9vhs7
iLYXLKaQJYiVO1haDTnEVJ2Ol526+Q6CjQIl+gqJeVR9MVNfECiohOJFagLRNSXkhJ5YvALx0GTg
Brak0H9GakhiGAjRg3axpaZH1yO5SBRyAYNwJZVIE+zMm9nBONLjVEBPdXxjUla5lN2omJcGe8VA
GI5OxF+eDeF3qdc1fi+Frh+rUF+IcV1cGfOw74CZyfeFmR9JmGOZH3EgVhhda6yQNBk6pPFfWJ1y
FMieF0OwobgJfBj/J6SXrKIhC2S4iaVUHlAb8VCHgqWaidndxYEhYHl4Z5cVJVehdfw4K+khk5Ad
yrikOemvBZ+A3MNMTffaEmsYAGEGEizSIYFzm4phOaFnNn0HWJA7Db9ypedWsBKGdTcPbIk9OorT
3WJokXUhr4EORMtKdGg8YTdqwea03I0F9kXCkE7iWW6CTD7kpXeJwHTWnkRXcZUcxijIg+VowEMC
ZJmPUwnTBp2TqGu4/Ua/9L+EmMQXLXSIBP0hE49XS7Q1i8zEBl3vzDs1rvItncxY8Vm/UsJt78DK
UkH0xTdkolh2RljbX2hPc7QTcryvoAscEdrMsSs1l1uFyhqlQkF0Fh2o4MZEC0IImZiY8rPWJOsR
SFhkN0566jQ6sZLZ6SRaGmoTAsq8nuYI3W+zRVXgoT1pwh15CuPif3TxnORM3FV1jEHtAxMV0pSC
oUTxj4uxgR568HkUW4mZSMgdZk0M4bqcFcKUk4WhWqgaSOnFfZ9asOmrLISQyIlqeKdRRbWbEAMs
tbqdG/m98EcSdC3f7tU/ZqdlrvqcL2jGFaspE7mcdTtZ9FPIRT+yGIR2mOK+wSUmQa5HFr/db12T
LtLYQc4ZPEGfkl5AKCsHHbzOJJ3ShpH1f04ph/3NgKo7S7sitZZteWDi/9hNRRZ/JPerM9aVbIAE
uuBAAdB9YIdT2QTfnKBs/KzQyqxt74+o2gOVbnNHCkrKT1xJHKxVN2CaPGCtOoetY9XcrRCH5dHV
P+DsQfc/PhDvnmTNjXa8hV5mNoc5nfI325Q5vfKMkJRVu6cr7Tj9xVxJajDMhvakhG1M9yw6ALFH
B+A0Nke+zORbWYg3tgiowq4/0ijZpP3o87y7EhQ5GGvf83WYptH/qD7fZKagcoiDG+pGdLtajHA5
JVG9xvQqHM0QAydElnMdhNfdPm582KBpfyY30MdRaGAtJ1BFBVd7Y1YW1VXsIjdy1ndhJSyu3O5B
VObBkOLnWw5PkEZSgPgsGjUQbi9Z0jOKXUs88sjbI/YkfRcy5pxkEw4lAFOLXpbH5gq7WOF6Bjkv
H9ckvbVrpuG54um/WANTPtXZgTuNS8ekh5F7aCiIDLny7nDaQNd9eoXnKit3UnNb8MOjkwRpdX+J
O8uz4oX4t8yrKxL7uQxeYds1OQzUFcT7H0ABXbBSznHVHDjoHuh2gN4tZ2Ug9RJ073xsSMtvJ0M2
vtIR8R8Li10rmEqjqYp22nABnnl92ESxRa0pu0LLeiZD+pzq/dftprWEELMcVIwuOVECwsnGT7mw
BnjV/aTGlm+W5E8VMblMUxgFiT7H9l7Vn+3a2fv95po5sXoCK/n3AtTo+0cSDNtC1pSHd3TMMNBm
nEG7Hj809a8+xkmpzzkA6OyhVg/3d81iPg0SkDtLJTb6hEMfp086NQIpMuydjPuyPCjPiwupxA8U
bL4+DSSAc34qL33faSs7JB83IDvZz8dc+oGgnn8gwo6//zRp+GwPrnxJ8Evu7Y8UuazzT0soeO+z
pQTaKbJOkjur6WXc9TOn+WkIOWxsvyeRO01eAr9EVrKkQhs/Uqb79oHutqxNQq/2dK0vA9h6caKa
6QGnRF+gf/FXb1yr+z2i4pGITFNUkTWEF9DKOalZI4SubiljZEqnz+pDa29l7IDgK80trCmtxqoE
Wj6kBI/Lc8/tfYVx5LLpWANrLaWgteefnsepJ54HgJaxQLMDl8cUGCKffMB7cAHHaRmcXTM2kw8S
Mcvy4ueVb82ONRERP+1gLvbVxIjpKm8J2sGbzjMjcNsNS5JgOLxP49SKs3g0nIQuagCF5ThUZ6o2
VBB5KHU31YEkXcCIeE1NpPV3LszhomQ8DmB2jhZdNfN5LIEjXH02SptnPe6+NohhEvEcLqyXnVc6
xDmUy24nO6MXT9AXtjjir4stdww+gB86pu2NdZhcx5y0xQAKACPpGLthNd1IgNIiDQBPqSGjYjoi
nfahE2ZPT9l++t+j519pyHVpag+nrmyZwSfGw/6jopKvLH+wB3dbbOfOGuYo+9HT0hO3GRORqF+c
PuA+PfjwVh33EzCg/dS3MnLgwq1cCbWfn6rBJM/uSvW/0N039TR3K4N19OEwukMx9bxLIQDiQdGg
cLtAtvPzkX1FdJNvdTsiBpMyLgGS4u9kP88uhwmQzTLGwxNSiZ7T/nVBNy0stNMAqLVRQzxMMXV9
obRYNLXSWS3aVWQ4e09V+57px0y6RPDjafp8xG9YGmO3ajFu8IfYI3eP/QKm4mJiYmJJs0Z/U6NL
dJjvBbAjb09QW1q+FNvz/LuxknLeL5fbR3No1DS0p89271KcEAL6q88PiVg2EhvuYlGyv7XsYRzk
q3CbRSxy9oAmy8q7wPhEXEecLcFT2WIhGInEwGr9DLplb7AgqB3loklz06Dx0Rv7iKDdPL+sUDa3
nT1ajl7gJRpycUhM7dE0yMe2S/cvwGU5VXhHAwMtA1+SfhgKtgq7usGzxw2C7eysOA4FnkTn871d
acoUjmg9IYSZTP4d3T+GUSOFWk3GA7eK8PVWb/D1jgxaebFBbcyS/EyDIcw1n4In3vs0uB/Tj/3Y
AdJiPVHz3SLv25uaX1NB2lEavqUueR7jZyS7uUqTzYf0VbKOcT0G9YoCv8gUgN8dbHDYNSlBem+Y
CRwgwJ8S9CcMuLqsU/Q518QKk+BqG5+E6Bwde9UfHyVKzNpCUwCKMr2oudl+43aTGM2ovL6Jp/+f
ceO5FuWIYBOencpnstRre98BQUhs5uzemGZ/1d4n7EUmoZ58OTOV1efbtuMYZSpMu/kEMbQShVg3
xXjoDB3h+c0r0fQNN+0TSVmxU4q03fFprPd7PdcBvzwI01AvVKNQJbb2qKq9Bj242FzkQAFIzAP7
Od1gLR6bM55Q6EhFk2NUteLDkg7pUzKs0V9eNmuE36rp/U/6aZO/Yht0VF4pSgzYEH8xilcMT1FN
nDayvXs+uCW0BOv2yQMpGYvBafc+h3jvKOlP5xQZy7F6MEzLD/3lRjFT+Ie4PxHZcaTZkRbmRow9
CWqg9VhYPJUHJy0hPHNZCGEQjqj71iAsiJTI5BbvrZxmFtBqXnZTUABuTtYEzWWslScI0RC+Gdug
I1YGupaFIYqqpE6lrOh8LTg40j84puUG3tqzUbqI426QiOVpXuKqy0IdmKppMFvRbXVWedpDSP90
v7m9NsU2AeOZr1KcKXU8tT1uNcoLyFCYzpUBrn1Js7DNYD053Ted+6uDR1L2mOkSpeYPhV7MyZs1
sGlTT2aqrs2KhM3Jtl9fGAr8TEdDLXKLGGlfVczM27QdiJW9N4x8DD7ftZdaGBeCPQiBjAWYg20E
wyLNXanEAO9icFJeWr2zJJ/e0AGI5QNBnkWcX2wbIXkvqyLgbKy7QBw/+1nEbTiYkLhqwnQ6aUuU
Tc97StY+6/jY3bIjqZl/gtaCnBcd4VR6Jc/FLc/b7XqqXQyzJake86GN77MHozRcS9NNuExu/9cq
6LE3b+pIdRrBXJvXMyUXKc61mpM5uOXExxufpIu3Ndns/2jIws4JQziUUBiZ5pI2piU66NlzlqJ6
IV6G7Zgya3M13uuCQJUY3qrZQ825W+q8HPr1zMmTiUkQmMiXYT6T4S4+K/agCIM16/dmIsEkSiWg
YAzJJK0zz7wniTPwaS2wFrLScT+OgZK4qxFlJbIaEF6ALSuQPu7/6y0YeENoYLZrjdlUSJCMbp00
RkuHX2EZAyGJHkovS0g/cSiVeAlZy+JQY3WIPyjVjtm+7yJ0fwaicbvTD8PBPhadX1hPWKfoOBoY
oLAv9e3IwVTDBQ8ID8X+5C/SIxSXlsAFpTFpyM4zLset1EgQOjXuA+UKW7uUh9Bkuvr5j8p4WKBk
WwWmwAOIkXt9xigL4/UuWu+VF+8nkdNcxacgbw2CfQC5F3SFx3FTtju0OtGWTS/13cjQ13GWd4sB
vgt+1mdJRMvPvJogKvLTDxX6EWesADM0nKpNx0bgelrYQfA3wTOhgjd+EjST0fuDu+BIzGnJECK7
wnXYyPprD+GeHvZH8rP9KANAKLDAZ10Gs227xIb6nU9y+DVifVjUIrGeqp4Phr3V0tJGfMDiFqLv
qqPN+ZxjDtkTDmvFfxPAlh6PvItcEFXq0Y7RhH/OhljfHcMJE7zZ2ceVdk/E7G4hL8AFYjB2B+C3
a4zEjD5e0xZUeAXEZGALdzI2UqU95/lY9na2ZsG11nFKhuICjpyDdTQJTj3bA2txXMJEv5aHhOzz
2BXwwjgqZjX/Y6w8UQYnROAQG0MmyiXYtz6CxP/oiOTPKwbChVwm9GNkxKcxWGPmrXaJSSBXhh4W
yJKnaT9sx0/TSuiC3VoOywfAk38DW69eFc2VmRYUzj8oAkfM68mOiHggti0ndL/eI8PXItl35mzy
emY0HIkebqt4oWSq/0/EydXkM+ENqcafbqLE14lRMhH/48ZVLkzNwR6AJFNBFrIMB8E9hxW0sYVx
66rz9KyKEyER/x7g9YweADuFxifNLi085fNWscHvvmEIXS9nRIucdX6kErax+yrgKtzqrmLMFA+G
xjQfMCyvGR9woKDn+43Sv8js3D3pzAd6crlw9qY8l/8UdK4aelqnCmGHkSOrAiXnKfEmhcV/zlxh
Z9WJrh9o8Ac5NewLA4Y5k5xWdJNLMtwdFvDKXA5VMXX3Z2IfeNOoh/x8aXAQULu5ugWK+k1Qi2Hz
TeHpjf4YT4gUMuNiqN6UWmaaQ0+1IMIm9NLD0EEaz7eCCeGt8hxPIE3XiyccdKtcqzawJLDKV8bB
Hq9qYzisWKkQOVdOZwRypptdetg2f8NNLO4zgFoVtIli44EAb9s8NbDZyCh32vQjfiBIwa6pBM7S
yt5su1Fdyi3D0+Z5nCMp8vtkamu8aqR4e8bDc/bTWT2RSyqN9re5ty3ZfUzD8iLgIOGrz8UmljnH
DTls+9Q1+NQJPv4b2KmfKnWe2GK4lrt7qnZLIY6hMl/ByhH3XWF8dlEPD23cKRk50sjp2Zkb9e4J
lpxohJA1QgxeoqvVbrycq4G2h1QnkRXkIViAG7l7jiftMgrXI3MQsa4r0dZLIsFjauUZKievh1GT
M5W8JyQwn2k24TLNFengowRFcm9qXVI9Z00c/tY7t6xfx+aueUGoXyqwMOid1q6YvOr6nMys//dY
JQn0e9tmQ5cCmKgbFGVkMTuLdzALZldiPUPQpCSz5mjOMQOgvBQbOz/H4WAJJCTTfzcDbcJIe7d8
TXB/alQsvgJvsd6fOZrmuiO+VHeoOjZ3xhclFmmhaT9yI68In3PTd9lReEfSpoKGGZWfOliN2HoW
kiHZ6KTYETHZANz0vxAI73ubTrI0iGL6gmbrcSiMRTcLwhZ3GpHCk6YZsC+sv0Cx4vIg8E9AMcBM
i1ru0cxyxDeezRl9BTOZZkGy0XzgKX7qkRF7cwjPOsDc/tER451JZz+mp/rTzLN6GuhHcqW3JIDr
zSAys9UgaXs8uevby3IAhJ1787dJfI30/oKLgd0cgm5d2Tkaxu+C0AqdXCLbrs4mXltqklMKCdFE
D6KHasWr+Bpr4h7hr5F2qSukjQKDnwKEUlsUcwt0+3lbc3QS0Q6tRhJOcPjIVKi9UQdTneEejS4D
fNfdGiK5A5XDiT16Mg7ymcPhcyjGz7+690pXTfTyPhnMUpCFNQTUtzG79La/lbAeI8zoHIB8RNlu
sqHDTBIwYVqBiaQj+JVt2k1CI6oMybaM5QEDaRkUUznxltalVy5H1vuksHWwUZrU5QNEPaWpV7rY
Z1qXTjXLT8kQ9luG7iqetYjtWJyyeWD4LF23Q83r/6CCJB/59Ts1mW9EgLXrjLd+0ZAonuMlAbuK
GGW9oxN1QNnsWRVdpADAPOakPdzZJbDIY115VG0gBqHqS8RKVmjUHJHzzJXYv7y3Fe0wwJRnEx5Q
CvNXjOgDDn4W2Bc6/9jwNMB7JqpmHhT/dS61g1hTEpQPdfQ2UPCa3BO9UT93GIPbtuIxII+XtJ3U
3XDXygWWkQnbDt0VHrg3to2OsqF0IVIq9V/4TLEm+DrN7OSX3U+UcYkihCxjjy95KEYLgOAy/3KA
9HLqAJM6ydyTW115EU8B4NOhlcXltTnTXp89y/Bj5VK9UmTl1CZKActYVw9Zvfa+K93/9xjypF6M
LEBxn2E1lcSCWMD+TPMIK8SFovUjM1edgbGSUv6HeUV0XacZMf+zc93kmJgqL+P8PV23WS9kWIWO
5SwWditH9hRtAtpuJltrydULVKbGVBnDYjh3oj7Lnb5f6yVHANQB0+ZjZZMOSNGTcIXzlkStXS0F
BPh7v5pvYi6/ESpGRbbHAgtibjcpQ5iaJEEkUwP5JzPg/KOzPuHgBU4Avy7BWKgArtjxNRZYQ48s
DpaDFVov4cgy4nSuQVMnZzp6jvwj00jReHlGcTtXK1RN8YzJLTRBGTnvCjKP405FKZbnzQx4cEO+
UVHISXTph73oiaZXWjN43hxKRbp8CzN+SC514c8WLV1FTC92X1iSGpai8//S/6LkjDiLrWmzo42g
smccinn5lyYeQWyWVoKLv8BgNMGMOSGyeAgoYp2oLP3EpbFOMzbohjbv4fev83xsdzW3lG14hwqf
5vhBih6oYrV3pBcxcw8UvTUFLn/c45TpFXOrFTyMx3h9+7w95GC37LjGjS5Xjdnf3noHJHgAACiv
KZVo7AYQwFIiOj+8YZFSfVFmqAE5/fk+s52UF5pr3W5YPkQaxAjSuJLoRLpSFPPgl1vUF0KXvjt3
qXOxQOSbdRVV+gDThRxm1ujBIacFrFBcXSkOyk/u/qMMhwME5zV9XymzSksyhJgrigjVpNuoMz4A
ZtW3M7/bDXTPZrOLxnFjqPLWsgQ1gq5mM11g7lg8MHtPJSxt/XayuKmxJsb+OTu7TOVTYHSON/54
ehCVvdVqUpC16wLzwTgHfESpcK9aFNqGiJkZbUjAvLZT4ro8bWwxqa9hwzQughCivjt6TDTBeJRU
A3jcKvJeCpnZMI947CmXcvj9nYZcDwnzkhFhPR8GJZGhNwl+hqAODFDvzuZ35Mw9uELTMtp3MOpk
TeOeUEJTOxdY2hCr/I0EOOlx4yom3ebsKG9SXMQzTd/HAO/Qcc9Vb738hkxRD5Bjb9MD9L/X9mZ+
hj2ugHha3MEFvG7Mr/fv4qadYrjTkyMnYxMG2bNl12Ifv7g/aGyqsLxzKpiEAe9Fu+S5s4BPv93M
fojBiE1HHD0yE8Fr5fjLFNWcJzw0IIMUKBArdJHvflrZmhiAncXW+A+Y6bmv2Svyai9dKMpzzZeV
sl5YLbOWfl3/+17anRWkrVOBZ5wM3hYqpE8Q3qFcfhldKyiE7YT8tzYiZuQi0xuiVOI1XcTdxIRZ
P6Nx1QUaYOCH3RhLtVNznDdcuO+hKJfiVmWfr443XLzFU4K7IcNTmcPY0aB9/QxrTWFA1013Iirc
4bd3UU128KMQv6vUQLY90x2BJdI6542eXEm3ZhsvNSzhGKpZZPL63pbSYPJVaJSK7md2Z+bjFEoG
5tw419RiCUrSDhxCJi33ExPvlEGw2stdEC+ubjU8RbWCFryLZ4UTdk2BLILzTDwBM73uugW4KdCo
JPLSz/C+iVwkigq7aFhZ+jro3AFVNzLLbgsYV9eQQwcmxWD2uqLpLwH/S+riWlBKjzxIjycMkoQ6
0y80JoleK7Mn0PtyiIEb8wk8ktnClaHPmGw7OoVK7notSsE4DlANVrU6alw1E4Mdvqa1JNT8Pe2N
N/Q+QOs726+cWVK8TwKGcuV2WNhBuo+AmTdgPGALHr1C572nRdnijjj7qLXnFwVL2larB7sjnhTQ
Sa2HqSAgILg6CwO6zK9uzQYRq/RNh9THZXiuf/tAVRUKVHsojAzmUhSGVFudCwkdplOntasD5l5j
yCkoOAOswaY2WTPOM235enAxkUf22P6j/div9PcV9zFUkLHRTUHRIobRSDel7VHEAD13lVPER4iT
5YB/nzI1UUuuGuAuMwKW6AGHx4l2jppYC5jsg4ZtL6UfVaFXrOlBCmZmzlxbPCVOXCPozr5U4VhX
KBqe1nQYTyLARM74Y0baxR0+Sphe1nRHtK7Ujb+MX8IiMSFmCFpHMeKQqlb0+l+VRZkXH5dQXy15
67vK/tUFBiI4DNlA+n2j+Q38PvnCshaYgTfDoe7O1xM4l/AcdlHXMc2X0jI9/SABAYKhfE+pCa3Q
RsSK1qxTVmuDcVp+ITuImB2iIBZ19tqtYCJsCEUMJ4YJd3ANSDzNsrM2i7ZzuHb0KSm8CjjPJAcQ
+9QPEICCLelbdSDbAq6+x4JE8FfKeLhTl9i7BW9H6lvsiQcWYezKfiGvSDgT/vD7fd+uSwUrGUWR
yzmAQncQuSbr77xka3jrlQPHdtarTrvRYQmuSZlRxUgc1JOM6h3vRyT6g1POEkDHfj1ojbvKqwSm
pbM9klEP2AZvD7zhQ0hJAeC+7VijPHVdwLLjCLEtmdFFpdD72ABzyTdX8vTPEErCELdxYQsQerjP
6ABYDQ/h6769JZVoSPNLY9wXoudtheeGfgtnfxscLbLKqe0cZvQ+C8PQkQvX1tnuGMv2PjLkR56h
wNyBeZDKbSXbLlR5Bnb1EFxkKXnIOIigAy2t2i1mjMV0aY4pwMjFEgG/VyWi29SPmtqqMvbteovI
5kgw25us7v8hqPk2knmVp/BFQVgMrxxNeCDLUuPB7zmXJzmRV3EVG6P6UW2TZKiCJp+SwLs+r8rn
uVsXaIrumwLvczdeddqADP0BcDSIvV7OYNP2dt8fb8DNMH+s2iC5JcR0T7wDDdLFYw3uQ5Yh9YON
56d2lC+FIYOeg1YEq9Tmnjk9pe10BheZDjHwm5dwQWyVJu+YTeybqP6+eVfHlP8abMBeSxE/MBLY
uSbW+8fdz/Tyr1TsFhGPEOrNOeWVUx4ja9SMobeMAz89OMiDhS+H+eaKCm3czQEXY/UrhFXYO4dL
T+ioJiEtRDa0VRa5mUzHhAUEt8Zk0FWMi2yHVezTLU8ogV6jQgjTEqTnExUEA41XHQrr4pV1X00l
pArJ/Q8DoqUZ2WXSczil5Sqo+Ch7HxSXNHHnoK8IFtVJEA2+mfH4oKS9FLT7r5DPzPOOjmcF7M1F
PwCgyfsJ58h/f859M1gJBMk3oBlZ+goAzt6fIdVmuSXRceov7mg+5+cY2YZGxfktYKOm43hobOt2
PRq5swwEHBxSaTxjvilE+nDRF9b0hS/sj0N7bpboXdlZbMHgedsvDKzPiI2Qql6vfYr8JYUNG40E
ebHSUr8WkRWm9mvt34W6yVXPSlX9KT+8kBrUu9E2dH+yIxhK+9RLheqDV+fNQ3Pe+q4EXz+cnW4X
TutIWuYAyChKs4yBLK30lTgy90am3Y+APa7Ik4Uulj4ZEjRQcHqC3fvl1vHEYH66PPKRoJ7/e4Qv
JTWxvpue8Ep1SbbSTmR+BCYRGTGknRIVW40pks+2+jzKPD8Kr4dtFZrC0rMUp6uYTUruPOIMObMb
+mXOMdcuADuoLe+SNrqyZFr3sMmhzGE1UHDASvxETnoTxhU8m3rvrwCCHEjeO9Czwb0ERkRdpt2D
yNkS3lrLBGpBBcq3TpXnD9tXmUtwAqhunp67TrKxwhNVXR/M9gW48IpB9qvDm266ypPap/kRB6oH
fgKSNQb4zJJvemgjU/bKO7nO0+f+yi0IXl/D04NXGcpCYx6xPdPqgEejJUXmXCUwRkCEMoiJoHOB
7zLCuRqkymJfcPPH9eUFaB8dbQFmg/EzS7w3673O7LfkJh+1yVMHqctqSN9a6fZCuBnXxQ2xXjwg
o/4HaoTxi8SLVYBx7isAjP66JPS6LF8uWftsXTkc8UGQFKIfp1dSCwDYTVDi/2qrXoWR+mQpA0Uj
t5WIAJ+CypV/GRJ4W9HZol457rKjcENzYUhmcEjvy8nd1DOE4JvdgOfA2QqPZA67J0UnTtAxZ4Yb
+tMvnVbx9CRNIsRMFNBY3QKLI4/zElqYGtOgkRRq9jEJX+EPM0Cz0OeECPBJZ739ZLqxt+KFAmsk
try6RsgOyYtmS841hoGY/uMmGu9mVaKR7GgW+h3GoWejGx27oecnScNFA+F63h3UOHmFTpRMsSsJ
o6unKLFzNrgCLAcp/7U+NPB8woqCskJH+CtIz81u/gmTMQOFtB8ZVPpOmTzmDZVRh05wjAU77G4K
OfHt/hrhnjhI8l6nglHHmvKDXx45lBfxgzArtIJEfiZz2i0QOnqT8UaYNFoEaBla6ozY1rl2rUQw
QiHz5X/ZxZ/lod+Xku9Mp6cpIAK2Rw9rRdoYHNmdemufd6XOG6SjsKDYiIjY5bFocaAvn+RhhXex
Hn7jQvN4I5tQL/6Um4iGjHXVyw6UNBRyVuZyG8szOJgJ/hhknMSGfCgoRPbRDPVeZuw2M4DWHfCn
UHcsWoJleYoVlKmfn4ts4UuiOp62nJUmu94gaafyZXjtJVR2Y6WxAeu1wpVIQPVWROmSIKY7xQqr
IfJShlqX0VOL5hht+mEvt/Uqt14StgpjoN+4FEbmGCc5bFLD6zkg8tm+/Xdn74YWDZyra/HZ3ZZW
Wl9/CuRLnJiOcXZ0HgchDdQ9G3GJWgCdNFEBgBHjyd8bEczAs+E1TSBjM0BNZtCMjfgvRqZ+dGil
tHCEGBr4JZgiJQWAg7CRk7Z2bd8/mxGWm3jn72HWMosyBds6Xh7+25+Nkuonn8RGMGeBFm+05lGI
UV0Mn9enPtBPCjeHw7xaQ1HqSeLgtht606T8v6luCzs0wZ5nkbuxSNVp+Rbe31ieS49zseY9CX1X
KM5pcOOidIDhlJbTA4iSt3Qq9DTm9hRkRXsLjs7DBVTlL79jfu7nawz/jYmckc0Wu2FQeZSs9gcE
jtT1bJcjG1hE8pMl5zrFQ7ezSBa8mA1gs0lFDTlc9lXP73LM8HC091vmxX8afmDugXepZFipqjbd
MQp2ShIDRBeIbUloYZXxDKmbRYTQIsZXdOoYgk20FXF2RLkCmCvY2i5SDakuMDOK8HYyF/v/c6TE
FqbaepWEXSJnjkKc5gkMjMQvDBhU5WOk4vNXvZPDCT1wEothUhOTrNB9rjs08z6Ml6vuacrBJBmg
p0+D6jvIccHWCQeUrfJdP0ddWcHXf252mmJTciUh3VpnXA6x7sfhDoc92GapneV/zuWmh29j4zzm
/JW7sRM0vFDaUVRcARMuTEuLh7PxhcrHf3gL0m1Dvo27oVwsO1/GsclS8tqJG1uzbSPPVRMaE9Kr
qDdmLeta0qFrD/AHWHYBjV75Yhrc6YxepdE3I5nRhiTjmji+NvILMmLFfqhjeQjB1LrpFSW0KQLL
ni+v/9SDi1JJPX/vbrmxdSKd5H9cC9WT6+2BOPqlkxxUW3B9vzgAkgdVb9lVZdPlTP7w+izvHfcY
30DaBqd2myMUfVBL9oI8O3xkktUe+IRmLMcCk0gGnlpQquXkH4jpGpShWJyBWHzlVUzXbzaYkThU
dw+vh5GFn3eXZfKWnYAlwd8dvRUrJq79dxJE9cjISLJ8INKzPQNKguePtxmBinE9nJnlyenF7s/r
e3mQwbK4iuLnwZYplPwNz3cATWdipZ1QBHMUJ2FhSOb/VfzfYHVQRuJ1W/u+fKqQLc97KF5O2c77
dlxpTfce5b91wMbbc25SZ7yM1ROY+Y+UuJqM8BPSgEFAfRPj/f6AddeTANSMuxYbKHL2ymBDkfP6
Rq3pAZat9nG4jVZqnmQ+fCuGDT0uG1ggqvvcVmqyHytJSoLtxDs6DmFZz3Lx4s8Wh5nxY3uVMfNa
yzZm7DBq0rk3fZeywY+xDgroj9N5GvWfPQmeFv5hKUm+zk1xTPRtYreHcopMGSWlE4NxO5Y2S4nK
d5iYdo5yiqRisgALw8b8wMCP0J67jMN7K8f/LMMesrUiP71Tz1vTYR42h97ujvLfIQ/iRoC/3fK2
r8arxKrI00eGP7+VNFCj00dkGFx+fvv+Sxw7tp7rcUxJRToZ0fsli/KICv76hdiqo9x+oJgG1DTj
JvRJOkAPQu3abUlqpEby7yutZGVaz5u5CGhIxEEPttNVnhKujoBX1aRNaxoxCaL53P2CMmY8cNEl
Jy9Q99glqiNWzcrhyjD85ef1UiL0Y1gWStR9rgY26TokcmDpSiw5IeG8MHGYrDfOLMghBCmm5Na0
cbIuxQuUwl21CLxYnHmq12Inz9ryxEZVqBqRvPfsURP/6I4HdogRaa+/PNstAj1clmEU2A0u8Iss
mh/13jghr/x14SYbTSqjzVoVlZV0F/h989TgzZiemy0jvwIUieMZNRdanZG/xs9yCvt0/ge1V1bn
ThUqjeFr9n07A84h3V5QiZ5P/bamgu+U1Pk9lRHsbPod3BI9SBZWUlo8JpSDCPW13euH+zhpyGn6
OvLg0LuftsMY+/arlB2wsL4badgBJhEMgTCvOrwCMYq0XXBuDfsmrdsOnFk7GOLN77k0bAnFxOFu
XdYNfhHp3h01cwuRDqoAjr/4VLYPLA262hvkq4WBs/228Us2GUZYW7iLEqlYmllyy+3+benyKyhc
5UNqvNxHAG4kBvj4LqJY5yCawwYqXVOpvfbsSc6llc+axlCYcxN36tQsJvd8Gjvwah7IpPbKDre7
/egohGQMkvcI3TA1brgiuIj9J4/nuptE23fVVXI1cbASRqW/xZoOsO7PopvjAhlKynVk2lgxUQCV
mea0pbJjVQtVlvLD3rNwD37YqzfOWZgGctzNqayTucG8muVevkrw0RYBQGOjGKHLJ/hVN9ulMDsv
fkY01N/7wUC3jekZ0DHn0l4pJpKQWuuJkMmGtPhc//W6xDszv+0rXMxbAeMoWTYFivR+x5xajrQ2
4qi0XsqnDMTpkEpdPF9JHd7quXoaoLbbzWc4yyOsnh+0nStAwrh5BJN8jrnpWzE8LXhuZpmkXPZJ
hmcNjRlrYrHs97PLtKCnOwQ5gV+PFOcH1Kod8nTZ1tm2VzdBpNDfE+3PqF5FdB27GJmBLAyD6TXS
6Bo9qMGVnJoSQm946hvHHhjjNtxl5MHjK9iWlyPeHdPo+M1Kw1v2TMcXQO5tWvZmWEvJ3J0ezWXW
OhUflBCWmO9Gjr4rwKzp74WIXLH6q9PuT+g/X7h6z91p3a8PHKDc6GwBgnxT51zfK6+dZyMl5tUE
6LP6GyNgVBeG/RVZZADIsPiSjlaimGjMQvb1U7v8IVaVv+H7qSlo59XECsy/ew6zD93TNm++/iLM
BgAc1rVNEcHKQA4pGszi8nlDmjQzQK2diJIGE4nKvOCpnaQwdOUIh64OAq6HUdS7KGr3wtVYViMq
16+I0s8qIgrkSoq6b5uhOzctc+15lHPWn9CAZdui2+vfOdkKYqAxGhq8AGFb3iV17g4ETzgf6AI9
2/W/FxJ1nox4hIZdOOkWbZTWYKSW0ksSO0wQgZJ3mO90hYMg+dfFEA3THOd5h07G3/9TaEbyTEu6
yuayuXHr6xOjn4Hl/561r0dZp0nfS1RTcgEx9kzcF7bnS6zsrUPvRq4b7K3B0wTNtc+vtu8PzEAw
CtTHnpxnJiNaK6Grp7pyhBcPOT7SjJbZ3M9EcLjxX3J9mRl6ZeJzDSnoEJ1QJTJp4XW6eV9d7/u8
o1L6W4+nCua2oo+DPlLJRcDUrX504GtG+4sV48gbftYj9lafmHY3p3RFR77osn12MqWSJekYR3Ql
PqI0vX973L94dYoEgZ0ME2mEATMlkRHAs7n/V4OyO+HDqNRN7ttccNNNv8Un2ijxmgOsWdEF1o9h
yI2Wt3GOypYYLt0BRX0V3pcHrk9hnxtHmcy0dcVBvv8wG6S9latSPMyFZJbH+h+q5e8SGXFjjr/K
vLpYj2LFbD+3BWtJT2f3+IuoxpT1ICEpav52CXeiH8CC0On3fe5dwY5yNQJoz+oxtmKQD9n3QKsP
eKzrwFb8yNAS8nGKB2kVc2O9aCUSZLvnorohYltSedPZ5VR4+iLAtyo5ZOT+x4VeKV0LMA9RE5cI
o1FMpJ3YW1AYihp3S8603gSJlxBldhzkMWM1xZcHL/+RK3pg+5qh89mmypkA2brab1whEE1iJq8S
n3UXq2XkeW7DHTQz7lWETIb3tdm3T+SqfCwqDxM02fWlSeTdAkj8NmgUOipSpnZwQdts22CKPxNT
ZmJzC6CWzhYl1AGzkD5XIQNUxlDeZuEBB/a4SZ299CKN0HKxk8SVi+ujC6FdqM34IBgv4ea40IrY
z5oYCyl5vSVDxa+wKVNTTcL+W563Resa3PmbcvRCTqmWImvp+zPevVkD7folDHVaovf1rA9N5oTV
CYjbpxIFKylPvX6cGfROVWMgPWNJjGNmCWKLqKHuzHEPYhgeZzYMjNEfwOoGhoLTau4zoik2bYCF
tc1ayU9FK5svOhm8KpYQkdX2i/QH3/l57/yGToU8q5DrWzCgRCPB0UydmnxVOZSGWc6o17BQcHwv
rzvKXkVgmmMbLQzF6vzgPoBOxQ7wJH310x/VflewBuJ3ROMcr0fg1h0z5j1p3wIxaxuL5vF1GwR0
F6dbe2VFQNqjIYvQazaFIKG7LFZBiE7Hw/bVCKLlFHAfHd9myBeSvQTO+daPwhhpRo6dSMXGq3lD
W1hzgjTlG+GnJgIHPkZzL54UW9tU4+ywhnHBhUM/s7HlFYaToxkxsFP73NLXSNDGtkI1qvz3NX8E
9KkJEqkSqA8dpyTYo7HHLM7exXbTz+SWd+7hBNZjA9ACCX6u0SZzakx8pUjpJm1Xt6C1g8c0Sudb
2Fa+Ynh2qmeQwRDyWtVD8zWjxHVwPNDQjrTJcYA96V/b7BLOOxx+cwODKOM1Qu++B2d9m6XXt3c7
m0uCMbgrxI9PqJ0zT2ykfmxqYgZ3WjMJY4m/jeIBRjRaxXzdttFp4KtjmDC3JxBw4aMr/jjncBQA
YHyokxS7F8xt5kt5RBEKnzz+gKqDYhoI7d4PYdFLwn0wFdvIQzhm9f/1hxhX6dCIzC/WXyzI75VE
UlCZSBg9qhpTLflGezQYQTBsADNu8yOmx6QFz8uOkC2LW1QqrJw/+Vo4sSoNr3c2/zHAQouBh3iH
EW0dt3t5zMfjeZazQnNjBSKUwBWIdIVsW1ZVL/Ri3WaGvjE3DHlB/zHEEI4f6ay9riHQFF/XHc4r
SJYzzQAgIZ6TMPHRbL0ojRyiz5+1OHzayWX0Y4bfQbmvD3bcHjMQspmThaCtBOy5F+S5F8jYsFFP
ApwsD2zNKLh4XUzBj00B8MKuDvHfw79wB2d+j8voTNfH368JbYKicaPThOpMpHKEyuAf2k7fqyU5
DBZSe7tg+915saz43z/OHOyP0nD6Ov7awaWVp02s/VrOFl+HdJ2XRkQmDx+w/2fX13yGZwxFc5a0
L3VXwMbA2BY2+5gtbdch8ij7/hnDlZmLeKM7QyOzbHHd1JRRF2kVVGkJkOieY7A1uh7YUQ1Ru0Ew
H7HxM/+J3PTDDZmtSz7AUyhygzxxENNUDSumd9Iqdf3kf41GFjFiIQ1NJqjkHBxIrVuhk7V4oVmd
duwyShFDifO3GgkjUrkRkmye3fFBzHcds4ZxRHjsHXNBs8CAqWYcZMaQBrq+juN2FhQ9NMzioSIN
44DL7YDxnbdVN3FNc4GIozh0uybsMk3Qv4jBKi5tRXl0uI9kmQdpcvMSzuYVjpVgsQfxes163ea7
7ANRZKphpnFL0v3ksJHWUcWFx9hL655Wu5vw9K7wjBT+H0X+f8Bvz1HKcS1oASGRf4kxA9vrs1e9
gIplC99/lxW79Gji1kKgeFUyoVTyELF/dVE0llAs8FVT54nVr3sdQi2/C80Od5iiI2VHcW/jxLTx
VYIYVBtfe/TKHw9Oc+HjD2uxJ7u6scbj4KxvYBA2oD/PnDjY4nTMe8+ALmcxpPrDG6SWGatBZCKs
NDo/7G8d8eGH4yr6FiESUX6oDjgi+aGw7l22I3JS2mwuPX/f9POGvpkKFdxvZxuvYsjI/cRD3AJT
4xX7fLkeGK8EIkk3L01gyjiYnQ4zNtUNSWWHs5MVtOIF/9QnNz8rMo1p39Qw5gtvfG3fVyzjfEpn
plhTX1Lzbnamg75H6nrG8H+bCUlFhzdVPdWgznDhmMnRC1VmjGAq0eGqHXmkme/qjwe6gaRACrix
3yHloWb/uOv86r0eAgxzDCaI99RloiBsxALQ/feXYA+EvF0GLnq8TLveu0yktDqj9yvTe5gM077R
y+2IztVTA9ihyTDD8aAXckmNv/cBkCwdmOPVY+xOEVvFuq7mW954tr50AIYz9zqsV0gSN436/ceI
eJSK/Exp+/PbzyC7FHGEH+e1ul+i/khdhguF24at7q3ItgPPjCNH1jcYZGQBBs6QNxW8wqA3I6Hx
DmYjojmCdFjxS1SqY4ilFTGuTp0deqHP41f0ZfCJv7ssC9KPdi41jjWD41XFHvsAYl5QB4Tdnks3
0MXjC+4seYo11I5tTyObnRz43PaI2cZTyXnjvPWmKgcYLUYnjjN8oQ7s1lmG/g1uQL5lZCG9gsrc
AVesNh4vYwBas52hZc22Ctn0ekOY6Nww1iMwGfoVaJFxEjZV/xpR4jvkxFSXeDhFnklBGIL9rUN4
QkS9CrZI6E3PfMn70unassolVuWITp+ogZ4p+JQjfsZ08uQh8+589ZCB8JXV/++JkbkWCj2nS062
/jH0TqtQcZ7WEv20lz/Mmc81270bqdmK0RTvWkvOACmC6/qRgDgU7iGRGH8Ko7w/yRvjYHP3AX3O
dUGKCtv7wGN4ruYLPOHPT5E2y5xUsh1O2PDAClafTIhm/br0D4Fdqw0FpwDL47p9lYS2nScPTBR4
bKEOv1/KsyCUn2cRs7Wmgl6k+cg5bgBTKaULTq79//wE81eYOCTcmtlLOaWXueuOJtAYAjUCyWPJ
ZXId1h2IQGPtLJhUZDlTzLDuMXbWquImx7mtgTNIptZz61Oqna2ylWiYmVJN5n6VpPmYgReBUS6O
Ft9Kb0Cy25JXtSZEAi1kIfekSjyunSOczPjn8H8J55X/u/dc0XnJ8KVWxLodjGMAjcU9vmsyJX2D
94WcYkvshEI1TDPO28suK6/cehgbrd4tM41pqILVh/YgyVuKZo5fIkIvXCV9GGA6ywkra3P7V0ez
8sKAvQHabAHjNsxUwDTp6dGEGBHxIBnF+xyuClZcm/eKnkFjCwiIlNTOoffwysP0qKwbPJFsWw+O
cK3plC1lS/up06f62VTj/WJZI4dX1/lJfLcCnFcLMTksdiwoYb1V+RkdQeG4Nx3w423G8Vlz0k5m
kKcfjW6D6jb0sh1CLD6QSsiJQNb6+ekqtG/7FCk99ddebeoiHu6bGmMAHXAvH8a4b/1DocuLdWzh
2TiaEDUWQVZxEyi03QO3KPakoCDyECEZGEanUeEvfOjXc8rOngypwsWXDo5sRUnfqevimnZvhwPA
A/hSTWIWb4XCWc3zeIsFM88NQbpaVaLXMOaIy8MiCBPUUuJLuiO9WtW59Y64tPxltG4HU9sgdCuR
MICNCbG1cajsMAPEYqRR5wU8LL6rJXdieUjewzBhG837jTKVH0SIG1G6F9UqyV4D9+g93Dsy1oQM
M+Sk0djpSmR4Yq57HZCU3GJfYmXhkdVAetMPt3xpyQUVI3+ZW+W0Gy7A8m+VRzRqghJm9yrgoP9w
tAK8dRBE8hYadOQX9WZ8n3gFb84McA60L9nIaDCubs0SJY03JfGePwuVZvjvC9JDRbtmWAE9OWiA
A7vrQGJCWyxtL4yNOHAH23RohkcKwydXqXbDL/xaYQ6z6HpNzNytCfny3qFPOAAIn1kKQYfCvSwR
ejxIv84rkCAjLHfpDCJ8DyalCLNENA3apxWuxxLKI0xkza8WdmkmaYFg7hwjwD7/PZypRu7q/pqQ
HKWbjX6ljMwB+06BYGtVZPgIxvPkNFcCUg/WHiHX3d+koLLU7IEe5tSErTPYAPsNl34CUJM5Rin7
lj5zVHDWkRa4XLh64ljX9WkO7u1N+Kh005sYDb4TUrJvr+SX98RSbrtc66JL8d96mRVcdAKRVU2i
rqvN2Dr3ZA68q6mNYSBkA3PteGaFiGALO3K24kCmBOHN51+H7VYkT/dZdNMsjXDRoNdqNddb0KoE
XG9AHXRA+Ky/PxDGGlLICefNYwEIaNefW5oJnOPeyl5Tnh7MJQYwid1+Rf2qiOVUEG4mkglaNPVG
HjK2YnD6va8ofIXSKG0L4IyiZfeejQYaFSucIE6K66/tHUWQHvptUHd/TS4tIjZwEkpI2v7imnde
pnOWhb1UVYaWDu8g3I4bphkKW1e5a2CPZTZFPDaPlhf4WoSEdXqLZinWEtBy201MFUtUhaDvjev1
mUL2F12t9LgpPFOuT6QGYyw42ebB3K2a1i4LjDv++DP+sc+0U6PJgO4hsDJKGFZuPKEE8Y/vYWfZ
lYhKDR+Tv78Nngp3efB0wT4Q1XwYr1PCpxZxJ/dzfMJjprxX6jRA6jEWihlQp8osxttoeYRNYB/0
RSxPxyv+zi1BVLct/TB75f/KbMf+EuxrBgBpVcYAoX1AWsPLN+Pw6UFK1RQeqyO+IP5FJUN5z9CM
FHXvpHvGJCJa6fVp/kCZYGcJILml8FN4fh2D/9+66EXf478nN5G2VKK6FWiziZJj0NHIvlRD817K
KCUl/iZl2I4T2Q3xU584J9ZE+IpYcgZeYXeoWZmDC6Cc0DfdVT81gWxSKSYLABWfxFBN7O/qajVU
vmRGDCM+VWuT4TWc+OF88wq+GoCgqP6Hb1qoVZbdgsTu/0eHHuwXTqfxR99Yy56dlN9Yng0Mjhmu
/5BP4UBqxGFo+DoiNsLpxt56c06hd/CRCfwisTRegzLHj9CNHJCz5Dwn1ANlptIuWbHl13N3csKL
8+eIaPbk56jevieWoL1q30n8NshjLuZMe09XdREcv4Gvn6OLCUepC9tvDtwdntLvUqhvwRWFAV1m
VofRwSFqEIXt4kbavfrvkkSxJEBOXFYXEFdvIxBkAnWi+qy5L3u3/YVtyTYcezuWd3Ug4fVWDsNI
P4zoVtROGqL9vfe3in8LaPvmSkKnkGbmw7juHJjq0/NSz3o6UU593pjP+AiDvHhHZOvK5h3w2k/M
rRSKQIDoY+I4v9wrUsYBQTmAaE05G0e4ajZLVnd1BDvRIsJDLHSoitlAD3HlFJItkuj1m5CULha4
8KHgsGuPXVQeJcQYfqXIw83H86Q25kApncbnwICdXJ6mbhwR9ZweXJ/CfD3ZMxG+zBx/G4+3xnVK
SCYoIKwCJhfYfbhQW9vPT3Hb8XFXxTO2B+1VMmgO4PrPiqrOFc+RFlZTCHYFTzZRPjVW1lCkau4D
PWRfP8rmEI8UvQ7BlXFh279yy7LGciuvdOg7kCPmRj1qs6qWnozi+ghgE9vypAO0FOiRAzqbpPVY
vJsPIMh+37id80HidrFi3sKxdbE4LvwLXMyDIXwwmGBvNrHa//LHcbAqv9xjYZL/T15aRnD9mI47
jrSLuaYH5d1x1VSDW6nAm4Rn1pxECIFF13fm8ppAYmXgQWEp7sCAm+ih2TEJ4+bM4coFwf5S2fV1
T71Sb6P9SWWqdeBKy2KeB67nplDYb/ab3xQUg6yJEkrDzdald6YSLjb7e5s2EA1FAwl0GY9z/QjE
yiFRZpvEAMpbmg9OCXh+37PpK4qYxU+yaN+XWrJCc4wjDZ9dwZTIFdzme/fQZt/NPwwZ7s4eK7fg
z0fYQJskK8O/iCvMv58q4RL1h7em3S6NzW5LuEWspZtK9INAYrpj33yjS8EwcoewItesnIniwrFI
sTvuVq047ncGl9f3vLM/pHQZQHbpgpYTgx6MeAKM5EAcRZlUd5ne7o3JNMbdU3c7ilG9i6IMScgU
aZ31qRYep8/eDRc0DvF67ZBH82NC8k+hcMdbw4XvizeHX4Wognc5hg//3u62XTSsQ8YWZ6OjGAWC
EHjPfMOHDBPfbQOFVqV35VKULG1AMQunMgXlLSrsQr+J+qdZXXcwAFbxCxMgROOZE/8suT+mBn0T
sUkSrNopfy/frqn0uUSPcwIDKb7UYu92IZ4rImCGdn+lHDFgTwURdV54NKos8F9x+rdH3d9aB8rQ
p1CtDziYHwRrJqshwd9PD1uySVDmGghylGvrxDoykAz56OmDOt9K297DRhLHs8zrkufUEwZAAApy
FLf6nk469KmMeWFFXDIubGibWkAPjqzXy6RYK+ONzrYAYzUhela2qS33QoN6jJWtaMT6fxS9sV2Q
Qqb8bitB0WssifPWEjlLLDL4PTAqtrJTwSD+nhRBzxHnxLTCp9WirEiTcB8HS/G9Sczpu0+Hxwt4
FwI5gGTrc8VpfqTeOqqETgq7457UBBzwVYmevJewjGS2j2k29XJi5IUQvESbPhBfAIfk80ObZGpn
grHwxrKCRczppfvs1sNX7OL6WqLYnKxqliKRNA4lNnIwszPspDB87mwdu90vg+7m8XdiG1Oa5FUd
x0UBt0B3WsFy9Q18mfvhHswBjO0VcQd0IKCPsg8EFYIqZ8xKulMyNku5EzwtH9GxTZOGCgUGeRbh
jjqeN0p+ItbnVJK9psTKY5t8HDIvbXSeFgtUAQcmi65B/Z7aY0anQAHlGy7QI1eiQKYr5qCrnFq6
vWGyIaBjLB761qqia/4dZRgzhswiCwvPvL2GKV6qe4tEyXM5PcTgmQmQ62iHphYy/iws3V1hpUVg
yBZE0dlUizvjOFS0Ll5S3u7bb1oSxzEHkueT68Etu37SGrxEG0Zgvma4QWtPzKuGgcPJBHv2aj70
s492vojN4BbPHa86icjBMlZijN8AyEzVHwX6h2/IJTCUSeGUx/ZizINCxCWhQDLpgiqCxKRlHypM
y2/xUelmB2C/GXtvrHSZmtzBSBlGRufdnT0OPgdXNqcOuh9YyDHFoMAKSiKEStJeRUtayfUWoSaT
YmQGgIuZj3MOkQB7x5g+4/IoeSeChJWVazQcBTrGxNWzXQa2x/eBt7aJDGg69OMmYmTlLeKNyq+g
3ei2mR525Q0Na2cpX2v1AxG2BgZYdsBGnB2u+6OH7AYCQY2Ez1/kdTQveU8n+JvtykCvV2OwUY12
PWx1/eTKInU2O5+17jlj6sRmy1CtKGeqE5PTlUi+7QZVf8eFBtxQaxzNpRE/s3J3z/Eq1hPRtCWo
vrp12yaCbiqZQg2/htK68WF4oB2J5S0zjDUfTIxilmQc0A6Rxa4xHuDNvzae1+vRB4LuVsdQSNi5
8dTvrMLhrVdDEe1VI5CNo3K+whH5BCX1+M6h5MBdXaVxBEIxFq08GxQcFnbfO5yl2CHoaW30Y6gy
C2vgro+r/hQGa2D++oOmchbXEjb6kZS9SP5LsWXBrJZTHrQny9A6s8QligdwpYkGLfM9DEGNM8L8
i35zF+27HEW3w2PrOwmBGagC77pExLt2tLIxckx7N7s6A+aBn578AN+QuHvb27NSHj6RYFz4Pusa
pUkMVqDt4+LgRSU9aUrWoigsE0NfmK2bi1crQCSA4aNNpPOWJuzJBQHhHa0SkdzDFP/JwEz8GC/J
le6aFT2lnxJzjdO5Jr6ODo9F8l93NOQaSRzb+i1YWP+t1O5nhY1kSRHHlwJCNmJ/xQ2bnGMhpsFA
vGBYm7BdSnpmRDif5aSRJ2HLRvak0VxmIQmkcSq2zdYZvoqtWGrSvkJk9ZnEyTVh2TGYiauzifZY
XDISlORI6xTwurGBAJmYc8pIr7Pk6ZFAn0Vo2ESSiEZ5eOZeDGL+UX9CQb4yCcGPV1jr1pR/XCE7
rRBnA63XYxZbE7P5wDABvCf4s+dMAPhvuS723BdSmqB73S+1PTqgceoll5N4qZIUmpKgMdGJmFHE
R4NpycuHjJV1tkXiRGiU5Iy6BHdru8cZla/QuyFORgYMyCnI9K5M5zjddIfj2jb/qSK4ggFmrFsu
o5NxTAKPdeCVs+eu1q/lFE/kbQby1iabmc9o2UpDPDs7nKk6wxIEZRZD8uzCdbXP8gCMCYCmq5eo
HeVjJrZBWVyNLaO1/MBrMOj4d5g/mODOt8JywPHs93+OaahM0DSG/Uh2ueGiBJtSzkySvuR5Wrr9
VmSs2HNi9h8moqjiszLOvIfe145ERthACZyZyOPT/TeZcP2zEiha5NLzqHtvQYdCN2PJ4IDXiroV
3NwIv6DcfQ2aYhertoQg+zZnQEB0hlMqFAa97J+xi1hJDNxN5L7aNg/ZTuYxtL5stJINF63fvHcT
DUzrilzVAaMA5iV4fEoNHc8+kg4SRYXslhQTLkQ99u1wIIeoWW1M/8uCNRt46i0dv2gDcJRFOdsU
0SPqXxYNuI4iA2EAlo+dFNtAPevJRHFPLA/cQBbsgyMZhNspVRSvfkEF9tg2EB1AX8MJ23BGf1Rx
BCc6KHBmCyjx4twRdSCU60MafNDPhOHqSzd58UXR5h/3TitAHRIEzY51oTp/xVBWhdJsIiEx0+s1
2wFtghDdH2mIdVYNr89ko5HLhKI3smeGezDMQpeMq7tUotfSm5VNcHo1sphgbSpTzM+66PStGl7O
eLOxLI1oyuZ+3PRvbr3F2m7NgrJLMX0/vC7eFVpICTUWQ02NI8+ufcdXEdHAQJK/Y+8bBSd5oUmg
5H5Nb3BEJ5VXDKwRmWa2UEvbMivgxVUtObpyrvzXKqqvSqPOq88MBxpkUrVaCj0C4OVui+t2mqYU
UTgJSsDFuPZ08W7Ib19OWaLZxEpzo3QLcChFyixx7dp1nvSZ1tyXjqlI/KW3ClyplTYK6WKyvXhV
TodRYRk8qberIfl1TJbTVa8SZ/8Gx6lMbqfi6PdupuM2kzDusMjeDAZS1xaBFRwcIChZ5Q5Ph9IQ
X0L9u5edLCP0bsY3f+lBVOboVe2J3GbNwu1UMbrP2AN4qwdpkLzVsPFFvxKv1SNdP2QNi4GPD4Hr
R0iB2/TIMiyCAkgmnbsvptoKSiStj4XT3XVIYBJ7mxAFPKiea4gtsC6pA3E86Po2No6oyDO6SI4t
me7kNH7WuuSJam7zNpK/hR3Tf/L1PsR1yEP3AhxGJkGC143HVIlhcfQDoz2T4DMJDY0D22jKS+eK
i9FiQEBqxZFzJ7RR7JuwdfoQI6a1B2ygrBO18MdM6soiiHq5w/U/2KDc5TJUe9evr+sbNehUJvBu
49t6oSJKyJdGmdS6kCuDCEPx2BeZYAK7GgiUOND12dG9OOuGhdCiNQcLbaWQd9OxvrQS3njE3h73
k1Z3dIsyaZWS6SgfFCXabPgrTt/B8RVijCOx8OVvlNDJl2jnVDC8rAJN/QtZFOXlIkJYRmGV/GN6
s6KhjN2WuzZF8/lEbpXp/qZBabXJjSuF6w8XBXKSDCYb4do2LEuf+7KxyCmAydkzRcsn4m3Af63f
7oRoew/scGWupByj3KkW4lkeQQp0s1BcWRRk7QLDRlF0IBFNUTkuAdmvJqeLvL1EsgFk1lRsPZ6Z
WCLKpOQQiwjdTCbxV2UDhKtgeLZs52ColDmE5sHvk6oPZjM1B/+HKxU2JHEvHorjzZtWnQQb6pUI
youvMCt91MiLsbKEuIxRxkzPrhOikdw9bi0LNQE2DQBsTJTlGHMoi2HaLQH5PYiGVNMf8ldQjIsY
RXocVtwYmMI6iFu1auI+toHm5Q0IKotmNzyEm27qlVVKFu9WBhNZSmtqDzxlj3d+ydijwfymYBuI
aW9OY2U+Zl7LygUK+uZwQAvZVT5DwQka18/neU7vGvn/Ha2rYPPDFXqZHBrlRS+QIXU2iXuWv4Hy
TlSIm9dM+WvmFptx2YvnHQXzn0t5DBFrXCQsKm62r0I5QRH6MAcvzEb1PGAuSsPpBKiDFROW5ttT
B2sTtfp/GgFAsdFg7IIfxGc013JpedHxonp/u6ePb3GGsi8fSQxFf59VpiOJPOha8iMRvd0ptijL
+9K5LcnWkuAvPfyfm69P9j304QC8u6cw4/Ft1DSEwf4/WnENkaj0bl0Fq+r3sT7R3LPqHndi0PyB
Ovha75bww1NS+hlyGvxdD2i7VPPy/+G7RAwoIPAjJTYzKXABDMM7oOCsqG4LGVK0XNQjQr2W2V+D
FMZlHopK6Ezqm/AjAiLiTyxmZaf+Snzdzbq7wduxPylJQ7CJOvfMGdL+n7cMK3LpKSMvElRQ/i7y
IbqBKujWFTMmpMHxVJiV2rUgb/u9ahzN+tvi3yp2PZwn/o1HGYpCIU1aK/cT/l0kkkiO+H874gbo
ndHhEJCgX66alBA1bTJDoJnVQrODwolYPGEwPyf47VQKEPX5VbpLnZfScWpmQCDehOAuNRxkNvXH
55Hkv9S5zRBwnq0ngyYZHoZd7uduWgBbzxt7uMOxbp2KNsDcjy7aneh53FU2riuHIFRoyPX49z87
dQTBrq52p88DRyDGBUZjVAvgN58TVKEwKX5OiBjRFIXD3C8qTkUIEfWmdbPW0mQazUi8tm17iHp3
qBaF8KZgUGxE1FnH4Vbl8NRpBcTk9kx809906tv34/4TwF7TxEMxcav2m4OcoNTZmWSiynzYBjq5
dc3fzV0zq13rm8RCIEwhY1fdmuSK08CwsVYhfex1JvczZQdAUDFgaN7cg6fB++UNXC8K2sa+FE06
Ay6rtOmw5piVzmaQ/HHM4UvR3M/LO9hdiOOPFuGassUb1noQZ0jKat0SxOHaHmIJGYF3sjptQt74
51+Qk3fSoYCZzE2uQfygDNPsgjaY0BJEN8e8iKheXmKUPPBz+1gISH/N8bFwJqlIc02jZ3g4P+2Q
4c6lVDMFBELwnEalLKpaVORWKDuWUX2++D6p1roR8l36ptVP04gOE4DPWHxlaJBw5wrDYBBeNw8s
dPzyZIMirEBWfmpzeKnKtXSa5eQdqg/DHQs8oYcK74qvUTCAUU6tjgirofqek38lWYue+Lfl+R7s
nyv0cdKb8Sf3LKYrRTdwqKhzLErbUA8/erwR5UNvtBtefy98ip75aEwv/P/V1qHlNcHP8XRnmwlg
JOurFhVaFN1i8lNy/Y+Jro/IzwGlleBKaCcHnsriNQAVlEvaYYjicZldDg9dAiXSJnTpzS+8RnU8
90gAWqWzuA2TWTAHKDChxIlN3wMCbqqJ0I0ri1ydcARafVCpGKFXQM7DqX0sIRv4RCT4G2m4xhc8
dbAGjGgAE6upZ/GOoVEgs/ZjpJx0uc8T/9btSLMq95kMvSyro10Y+Fcbz3RZQ5Tgv0ZEhYOeNzo1
gdmLHEY2gcBB5eB1H69OwwLAgFOVANRTZtcko8PKWXFuVRqKX8MhWOM0x4HoxiiNGNQSv6qHrlA/
BqgjLluLIKuH5ivVwzqMQBSX3/7F1LZ9opf3ojz6d2s3g2qh2tLKfEpQ+4Cr3JS8foF5DFbvNLdI
LnYytskzFsbvExqf+LycIqJwoNmZdKQlTQS2tqf3YzUtJIarEcvlYUcNstcfA/T4uemx8QuDRc9x
KIgxDM47nwvZlf0DnZZWxLVS2lxTCRIiIZSqynK9CTFSDRCodVztppxjp8ps3L3nWRFrTVtVtE9d
4+h8r9IGfJ/5aVh1tUgJd+YYeK8slk1L9giZGzcDlojS+OiVXdbhEHsQma4jP18C1FBT3CA6ZBEY
UEajvQQiSx/A+OXIATGyAXQ+ZJdl8ncEgPLzXhf0cfl0GwyELMf+/WdVNWzmQRiarO/hysu3NmMP
sCxKrEiX7F+pVO7aQH9PY6PsdlDFEAbZkQCVE6IDM1XaTzGkXJYr2eBsWssUGY5k+W+7D7fbJoQS
F8IQUmJ2zka1mh9tdD0bxUEmMVZspTFpBUO+gl3+WAmTodDqd/6aQbCYPxHrX5t0ghC7lc2OJgp9
NzLGB18it19KOShUO73LsMzkUwIVk3tHDvQfJ8+5Qrw697ctqfbhkRkf4bymCSMIHazynN/QH/gO
iKxLQMfPUpywEBultsAOoX39d5VXsDJ06LLl6KNvq7W4QEg2jR/WdW3cRCgbU7ztGltSwIhbzgaS
vYW6RHQiVWLqQf9LD+YT+ykuFtW+EJ8RCFmUFxLYDBU7EldIQBehnb6B0KBK6sdFmDx6uRFrCSEQ
IF7z6uLXdzo8KmQbpAD1t0jYuUTiiMNb8J+JbIS9uxkf6nf30GRGxlb+NlbPwWgiPV4tf8lxQwGU
m04Sx1P/18ZyWi1/DpxYOXWXTZCT4TZNQ6ZIPlkRW8wM7VDGwOIHNbkP/KHU+Ar4abpDs+Ye/WLy
BPYKF7bPXz+VC2oYWpv55DDpeZW8M6lvAEcv3cqsJIdrThJw9vCetvdBjnlrjZCaEwRViFkj60xk
ub3JH7z0sWsLLt1vRPDi4f1MP626EKexRldqQOxnblXXy1YuajyEF1y9sj6uOp4hptX41Ohu16wZ
Bk0bBAhJzHgBYp0Lk41W6V7lI4WHCs7tVThEiiSDBcDpVOvQajLKrmDydVdYak+vEi5qYa0cHNhc
oiIt07Ql3Vubw/LfHmt0b/uAMnmqiymmC9vQj+92UNPPEC0Km8hEr/EkzdCOL2dRBIDJIcLouFP6
tpkRH02TQmuVGXA1/JJ77HZ8RpaY3A/UhrQm9+HHVM/Gr4UVq8qO2Ad6OEMrgSGZipo105OE2vf+
WU046ViYQ4d34ymT/9sPl8FC5CNRNp3TD0f20kqfFOlD6qrauuPKY652fyfkkmHlh1rF8Wbquh6Q
nqNWP4f5KeEBr53vlS65rUfKV/fJ9Pq/awZiQjLcQauMnz5qS9qihSasFR/3AK2L/lkE9DwOXmqb
33yqhRTnkMH7hOx5DWaISnRsleNhO09wqgSDXx9QE6L21cAcn/fTssW8CPu4ZB4s1yu71n6WUIWz
J/lmyyes82KPMVaQZO1uIG+7vRVE1A9PNKqE22XWP92Fg3qwK39xzOL+3mJ9W0ZhzmLpD1St4Ola
XvF+y7O4DP1Jd/FeeSmN0USN2cn0nJd14z5ryljadi32if6uY9iNKIfl421Ict8LGn0gWfeeZ7bX
8Hej8Sn9ogYJgSYom3Y+ZP6mqoSIf+5GAHjFuPNiiPCVNw18uoCyCfKj9bDXy8s8omDePbwHd8Y8
ClYwA7/Pb1kYpwjfLs9q0VpK67261HBJoj6tq/QhFZA4AMO5aiWmLfxYbuhNLPtzJXxDGXKPyDbM
NkLyRYGiYfTmefgsOpHFrcA0tTRj+3zFfFMH1nn43VOxV6e6aE689XrGQSGQGrh92k5TAcEcCmx5
ekBJexX+S7ajrQ7LrIDw+VxSl81diwateal1QtYMJHpDKgPc3lV/Itslj/ffGEHv4N911Z1RVnSf
zd2bi+Xj2/cPLVkLsuN5y6rXPYz+wLovjsLy1Bo9i650j85Z1X6CJqPdhWFNRX1T2Am0B8iytfa7
/lJg0d6h/s9KlExuN/LY5uHkliuXYdeQv1JIblCUHeHYy3x7Tk1fyLmt+Rpcamovrc8/12zq631E
b7p+xbywA42JJ8rORTVZI35b+d8KrZjsoTikgQU5NHMcXDTERjqchizgDaWyPpTufcTIbj7rVJ3n
WgROiiFCxxFndvC56nNLLXXRcpX1TD6Am5pUKCbapT+tVR7IVbXhdPUqO1t9NMmZG0DCJHM5kAvf
CJQTsEZRM/q/rWOBcRbfiUkznV4V4CyjdspOiFOo7K6cXuW8524CyWhDrBTE9JuS/yZJlVRLWxRv
AwfQDB9FnhxPbb/egFdyl47Lw7IjTSYB3rgYNAU/Zd4BZFmuy0QFFa7hLzXbD6Ou7cxbRsaEorMC
PL4PoE0qiW6xJ4+zDnc5BI6Sg18b/5syy6ektjGPdxXAVVEc2Q/6J4qeh5BwazsUxfUXBy8WyqwF
Ap5CUSgMCEu66L4FSiC3p6YzxCdD09Z0rFSHraA4i9tV4MT45zaavMDeE83eC/fdXcyqhmAETayP
gNAQj3rQ/hmW4Y4WfKYwVBekA+GHOEJYe4BRkFJnBncgIF5BnoPUq2+ZvGdq3fbFe71EYy3QGAiV
5jJxv2sD7UXUj8vETag8GYxbpOcN12F4bxItztZkH5suQchkE5tZFZdWsJ9hG94SDOYFIJ9I6Htn
EeZsJBBXhf/DPZiQdT5/xidGBHyEgPplgohGQYJXOdc6RjEgSqXuTtoXny3XOXld2B6Z7q4Zmyli
Ax7DjUz94CkSLxwqMdR4JG2A9LtJwytKMTGlnbw1hBTbRryEUrR3BnjOkVzMj32NnOk68aj1HMvb
iRWYffSr3WIcXLP8ZzfV5rRqRKenjEBqjsuvoBklhqAcKbyJc7s2ia+ApMcvU+WNI4VjVukd+va0
45CpJRdt1VnImtDT4fVe/sUyGQQSn+s2ztgvlUmuiW47Uf8aqobAcSGUxpjVeuRek1sYJVkSDkQh
rGf0Sps/BYy0gOZzuBI7OcXw5jIZzjXAq2jjx/VhodVw2S0tzyWJWQmibEEagwCvct7iFbK6B7WU
Fkad7cGjgJ2N6zm0l7kFxa/yUjEygmuvfS797oI36umgjGfv8y7ODjihHwPhJDiLpgUfzueM2i2c
XOyupOwafzC2MROmA3DNrjMVejrVO4axAlBE4d948ltRQTrFgy1RjwoQeTrv+EXPAAblaodL/ADm
gDV3MPc1qrZcbc6hGmMF1DGh/oM1Fy32e/rKpqVwkdXa39QsPrYBOhdLzAlDAZpoUG6ygqNbNJd8
wKw39R1IiYjZ9+zZtkzTs2SLemVwpLW3cqXGum0KHagybgdLfnqydlX4suK57KCupr0uKbR1wLvr
FxkTm0MuJvRlTxodjDNIzWImcsQDqLWf+Ns11QULFE6/50NPUkIALpdGaICvkxw9YxOKNmik6u4M
dK5/QOV9fCMcX50FDV7qTOYUQo0wYs5l2c6Uixj/NJWJZ29JEW6/ayKYdZQ0YP78TZyoPlqfQZJG
GiwAjicoG+ifpMSKCvfAWT8BCkzD6zfajnngUjogDRCRBoDhnNGkQhwLkIaTyBIjJEZxKPhqtK7X
c++T9oEI7DWDn9hOnXsnVMVcLRtrcUtlqgJ5oHaHimbq2MAM2UNZGQAkgzI3IDHHxl9qfgqQjTVS
0/1P25Y6fRlImz6Pj23Gx/7O6XZnVPjgFXa9TeIw7Xcx1Mw4CHijIMGtc4F7Vh+AdIM4QZqLmbke
BdyjCvahlKMYlV1a5T/PktfKVd1MtFfEOw0WuPtafnWmtmDAF7qlIg31zxuqtO4A5BoorgLCukfy
NzGIrwlhI5BO3XCfGr8OAsHHfzLaZcLCAbV1rm+Jwlf9srQvQEWdd+ObC/7UjNokUXcZT8pO0lNl
zEABN+Yslhuwv9jIN80RTyAiNVnPYBwE6e6u14ac2tZi12Ew8FLS8LLVnLe3Qu1mAm0UJlp8YNse
33RXElipPjA4KzEfbhX9jsRfP3hJ9UJZumafbvcO+HiS7lrQb26aFXycN6mYYVa4nKO5DQWyDXra
Y2ckcIc/9sDFUyuYux+ncV7iWRKRsQ7wk4DP10wQ2XqyZxxSm3U1PkrwqfZmCAa8FowhPPyW5+Qv
BQrh0wOdg1+SxwFN4+wrJaRDYKqsKyYt+85g9EQn8JfLiQXUhje9bs05RgHBfvtn/klOPaoQEneN
do3d9Md3hVYYfVcC1b4DRdYFbnCIncSHnMI0IBBffeAEevh2CGrwxn19s80m9jDFyLY7k65hRKp5
XqP2LmwxUyIk+2Mxpdb8uqWzckp68gXfLQbKrvG+Gcj2Nq2/yImIma6+3u5yPkkJMIXKM2OHQHn8
qtRWZd5uf08HPi3UXStyJPWHBQtcu++IIvrvPGufywie8/wj/uLFJXt7lexC2eEGGWP6wvgxR901
t2BHmGuvjodLox3251fntlLLLYAaNhoaUteKYaXgc8rDyqBXMaPOBhvNPMNv8WziDm74Dw7HU/EL
DlfI0EJCKj12vOXevsC1FMzo4J9tD23UkBqRNsToCPLH50U/sPmiGIzpMYljc+9BANSQSeap+8oL
wCOIVJOEq1ZVuqqHtyvhZEeYoStBLxEpht2Gw8ySEWPJCGhOoED+dtLPrPmsNmXuMeHgXH5DXjO4
kKxeI5AsxQP9+vcEQI/ZxE6U1p8CLTsos24aImZJnU3oRRpJvvMalKcNpPNYTxB2hZxmy1gPZkYI
ytip9Av7XPYFlgtR1dydWjf9eNd6nsu8jUkHc2j/szGJfu3jsj2tIBt+U2iGUH0/Vuo099xCRVV8
xgidZn207+IuaZhLlxYr2LbYYjVjiDNif9+kAAtJi2T3kD+W0WI+a5lxyCeQruccZpRKmLKNWRY9
++xmdcT0sJ6LjNARZ9lfqHPa7eGCCxwX7uhIQAlILKeW1MwrJ5w0EJ9fqmAEbcQ7V9Z+AcqzLdKB
vxSnlQx6yVGph/WYWMPqdX+XFTXf8p0TvXqPix/kNmfJkKwDacgdsZSPeUjjVhuKi5dxLUpwbIpT
5ynGgvVYD/ax+nRf7+Csq7dpEu82eZfa4Nki6jtUWKI6/ithitRlU00CF9Nf4qRX6cCLoG3/Dd2F
cTuOMSnCgWhuzQt3oCpNPZ5KDdpyS0GdpvqamCu3E/xWaFSgb0OX96XDBa+SVRQbo2OyX9D8+Fm5
TUK1Gy5+c3OBK9aRigAjZGSLLPvLRHqTPjInRK+XO+kXG9qrX9AHbnudBh4hhFYuf+EVKpTSjtV8
O99QItK/nydUu+403ugDGks+HRBPX0sA7YLlJ+BGpmkW7s+Zp70Dr7kfmNi+oGVVPFb0zDPUsKzF
aRDwlrxlF3YSy9iQyN01r8N0TOQFw+9M+FVUURrClK78JEe7Ha9YP6urLKJV6j/FdlankG0ddRyi
w5RNSvkM5LnzBb4WKJvhDcIkr+qUnv8JDqs1boCyiRLWyKZwdsEWNErzMIt9EmcoPIu4AzNPoRD5
jp4RuvtTsAPMvohM/ofz7ZsMKc6g75i+lok9al1xhSwjKE/x2y/z/SH6oL6lPQMuW4mALGgFsNHp
ysDTVJMEJg8sdr9vwBVK8nZEqLQhONEg71BlTfeDiuuEWbW9aqisrxK6kdXQdvgNEFE3XjNgBYW3
y6HvrccP1CGBwKhyl2/Job+Nwcxn2Kj4xCgB8sq26iMKhmryUIKxiZ8oqPchi2WMc/2GAHN/38LC
+WGiIkiK6Jw2N2m2EaXsWVHTMbUKu7AgXQM/RTHQP+tzEkPsC1UiX1dtSVMYKSlwhZM/4Hvb7zyK
iVUlqVnojDGtuaDTwEKLhC0ORkL10ytuvJOgMDwp75jrrXBkLFPS5eDzgD/veja5aF/D0Mcmc6ze
ddpA7wSZ7w5p2VetKs4BBJ7N1LoILFifgmBKxxehAECHFOn0whfSrx+bmMF2eWKqn3IVgbShbWRr
ZfQhVQ0vscMIC9gOU4h6JaRjc+zVzAE8kBxFInjU4ukZJFZ16DmvEw04F4Wfcj2zSF1A4TGiY2tD
T9o2ZCwkQEn64PdT0Mk0Rdi2utv9fwHv0p/NTKIPIOOgg2lhOEJVidN8iV/NX9PkFOMlAUzHITfa
drjkk3h4XtDFvQIOM+221SU4G1JduCY8KY2XZ9Qk1u7noj/RZCAiD/ESy/QugNJErxORbZraD4Bz
atXE/Or/RTh9Fy27qt3QClUU3/ADR54UoR0dZcSkCQnJ2KOkCTIHdUNM9r6i52+hbFPRQFXSjfxy
nu96N4gP+ynyZgNc0Gw37alyNDbelpz6p9vfXjv8YIGHdZqcEs36MQynkgWfkwIZwY00S23kfxEd
q/Fsf3MLpsAoQpHvItAhysF/9eZVQK6kQbRUQlH0DfvK8ufK1t+PB682VuZyqu7dlQ4uFZwsF1BK
L0efQ+VenSJx8c87Ko0jc82L2kOdNq36gFaxzn7sQv6Q9ZOGBybyMoEtyCtyUqR7VUIDg3F4cty8
2OsrBc58oqiFaMCThQZWVRaFd5Z+OR69Qy5iKJu3rQuNRtGwHBPcjagRIv77chMnRk9vb2mYoEtz
PZ5WGe3ZmniBbifGPtxHIzKfRsLhLIFh62NVvEAMGa+aMtK8ko020lr7KQm7RVvrBXvkmt+3q8kx
V0wxO7n2MaJlZkhvraXDmLREqTq5htS0qXBfp3KTUDbaIIdrsmKF3FdJ8y3HuVrIX/u98y00pkuS
lESBtmax9Ix9otz+JYES3v1A5zWsm9NWDSsrKMeFcWOFk0Fowcu1b++7kqhXjVjW2n7oDWTZSEK7
W73fUBNVHm6VtDh84OWdPvaFcRZyyP+xi0ARiEDLwtI3FF1yydY+ErpM8TL+MtIAe0S8txmPmvU9
7Gmtf1K0UhJlSBBUvon6qlN7kWxUXO/XLUqWxWu8QGIpHzQZAkxifL18RJ675VS3349JGeMXGenL
Z2HavVZ2KlpJCAhacnXQUKuWVAaqhBCV1FpliOZDh9C0WfTusuZf8lnIRx2jHGis/418pw1H6HVC
FB3xoJQTkjCVgFp2RbyVgeEelWwzYTYOcv/yz1I5s9UJXjcjgGibTKegAzxskMzbkpyrYfpAI7lh
llAtY4Lga0SOjeNDnZBSqAC87J9gz+jwbYpKSVeKIBoxNnnQhAv5bdBEUlSpy6kq7nWpzME0Dmlw
kPf2GWT1rH/eCtFPhb0J9qXzahuNxV3maCpyzqfHfCyH2mW392a5L/EvvoUNXemSBk7bJ4jKaurA
zfb8CzRxPGaRMznao493EAUZ2sd1ysmZV7D9Hjftzo5ZTeSi9ympPrExNn9HLtVVmPhgsD67s/XS
d/T97CfscemmDLToX2IVjxbF9PX2m5xONcjrc9lHzK6N4YYo0lUP4ChHh0BlNinZqot8CogzBM6c
nqBB5c3WQyMV0BQQP4MqUQWj31fpVzMG0SZCHTVkXU78g4MrAA2ys62ssoD7I/dQy4NTJB//nPZQ
xHcRi/50/Gw1n9kYwR1lXV3WINxd+2RABko+IYDLXfQQ1ER4ui0EOFkHZk96FDURDAPNrhOlRGK4
0atqdEsphgr9Awj4jJRDrpDGSXrr7crnW2utzI3JlegJNTqXFaTx4CAXnPYYj7edX9l6lH7lxzWK
w0nVNrR4EHIKFcg4eae4I3Sx0T7LA0g2olGejnGft5TKdyAlPfjkIB8oTZXt8kSYeI2+Ej8SELZF
wQKZn//S9Y0qjJA/8qMNBBVcamfK5vXPpWKqCRhftJLUyLRKcwAI6DvDMN/1hIJiH5hEfs+HMAcb
LuP02xiffDumCTvnE4JGjrUtB0SfuiCLXaRPxfYi0Cehv2Qb86/bUYCTYBDvlHxMLIcIjikzoc7l
CNGf1WXYHgrt1XAIqbaRu1SSau24coW2b5iRyVqejTGtdxZ3WyB71TWgyW+j7FRNMWU04zVc8PZL
ZMesbKRoQWrynTKX+VESc2F0RQ+8hUy+YW26JwXi5+RxUnzVau1jjKIsuh/zBqlPNGn2vwQLLJu/
jlf1MW+2kHWsSc7bVlUb5shh1JOnH85dlL0mtyz3RMKt21IgxSMCaVr6ESgPjRe167BrTdI6V+hb
1VzO72mr8M+PJvGfE/yqMobkCTO0wkF+ktfAskHohIXBiO8DpdlveoAyzLMNqOOOTKoMFVxBLuca
GjnL5iLnoUO8s+v4a5aOZwKwEzcKnxwZeJTPNveh4wwOyPaOw03S2NCUjXtF9o3FA6GVEnmLS1tB
qrFNE664B7yKGM8NA9EbuW+2Akt4+IZ9Etos3wwtx/9QpdxJ2IIqf6cm1Hm6Elco648B3o22dSW3
JfnX2BnEPf4wfZlnlpEstPN/ZhlEyeOMzs15rqP9y9LsQ0JaRSDoYe20trr68W83j+KzhvGuX5XH
nLTW/VWRGdIi2fJxwgl6BS1OLhxEHy17EPaUCc2FPaOD5mvtARRANcBOO2UYWmUTFAYcbShtTtQd
XKbvCI1gcKsJWV4DvkJUEFblsPGSJsIGVMa9g9zKslMYnixB78JhlTsClXPFdbN/pS5l6u2NFCv/
TjKWg+/ohTTA/jiQatDWU9XHlzkktBEdBnV2HZtFodTmhLxFvmUosg99VAL3Q/MuGGsG0XUTQ9Ur
G3xgvyY+Tj0gGYu5xPDHsIf3Iuf3Db1o97zPCVNwPvOAQ8jIMBhYwIEBQBfOS+AALk+Ev60e+DQM
GjOjtQiaF6ng3spj4OBG8257GSZDkXbzP1PzgNrwv05DK5zTIasFuCEmtnRYpaumm5rjRxF/sqXv
fCu/I+F6lvRCgARgO839L+V64KWp20n6Mhf5ACPweBCBnTByyTFJS36lCGXyD/3xOIfdMh7dI7KR
TUTEOVZEC44i7QJQG7F8q+2m2HDiEjSetnjUVs7kYV6tO3Ia8BlPhxhwIB8BasA+eJHOKuj3MGqj
gPg3iqrHIUffw1ykWrnm3EbuiBm8Eud9y64BgZs0aKL5AnIEi5ParAn8BEg5jG9o7d2DRr3/PytW
bWKira151qFE5Q8qZ4STLXiYzQTfiXlobijKhic1LGtyUG0om1JNIgIHjwUhYKzCtjRkfwDWFgIM
O4td+St2iwd4gDYVnxmN9M1xuOeTvvb0wqT9YDXSQy/oanh9di3/iu+NhUpNZqwNEOMrwOnXKREG
E6owBkA19KkdUCvh3zuUtqrosA9ASm9sZTPIiPpCDoV2qd9peIoauTXIOFUb1PBgkjPuOjc6O/l+
KLTRu38O46mbTXqLDVPcxA57vTjsocLYxKFVyOPf2SYarhMMZqm5AR5lv7u9O4YIk8PHRcIoYWEV
IYRWNu5hwhzw2N33AgjztZkNv4laVhGxTxoehoLMLbxGyVTMdv92cYsDg9YT9ZtLS8ducakZH1d6
dayVAPbNwl395jvT6mG9E+vTUzj1cslTRVFJSNhpAGS7JqtWsL8WtG+5oChYbcd1r5gkGgxDpt3s
02LaBMdmgsHJ4GRYEguHW/bpilBnDk/sAakog27IHFzQHtaNVdfIWrC4LZXsNuxWsjido7N/3VEJ
dIt1Rvdubb9qp8OswUB3gTEjGT+C5AL2IwDJgwbaKMWG1et9Q9Q9/qHoZxZoo8H3me77sMRZshJo
oJoriqi0O21YlGktZuwU1uvgjihLcepWP6CxrXKk79eU+A5URF7jM+8VDsbd/UKCuVyP2eRJlz+p
FiYdgSsV9esMMYqaCWCN+fY9wqPjBUNM+Ja8xCtiiWF02R51KI7sHAHp7bQkb8I1CIoUog4bwB89
DJY5bysgzWEDY5mv2h3UajEAxdOUWETY7woEmMjWCsTNHKxUPu5lT+X7vE8b2mXwcuVbFkgBMgUz
J5cQ+Cv5/q3UeyQkHoXdSZPqrlhkPg6Tu8kJYc2/bEn15Am1IZEpAgJrLDggDhLlLHZ9FHCVaGh0
MuJWDPg0psamlVbgbUY8xOL6QKhmj1h9KT3CS4i7Hp92oCNFITGXN2OZ8M+zc6sIzc77ncu6AITW
8UoA2u4jGEgGt0mDTzFqZ7T57zdgEd05UmsVz8xndpViNOsSVAv3b/JJWR84XBuZXlsiwRAG1dLt
WMqb4pRwqz1L2JIpy4R/uUVoc1TZSn9ycpxDs1SmytVRMz1GU8R1mAYqTUudte58qBdSHuJ+5vxF
hLohQ/Vsp04l4FK/cb8LnG46yWuAeWOrv32aoOJ7dU9+q7tGse1Ut8TYAuJ2gYjTo2qkkkFcQ/jj
nD6eM3iY5Kj+tbQMQ7WxOFsC7iF/PEiwvPntsF08TjUqPdsvAktKsr8LvaVH9unK5SXlu9aQ30Ir
sgr7B+OP7SGnbP/rpkDtHphlrTeW+qkvmAYe8qEWOjaZl5V2tDZCE3I1vAfzS3GUck0jcQn/Y+LY
AJMzuvz78OB5KlOz4IxGfyeDrypH+1Q9Alg/ErF8Yo8IhmXr8scRom8mkabJB2YagGjPK7GT/Y29
B6KSSUKllJUF3V8gzt5KcyPVuF8muA52sfPh6T0SkaH/Cz7LOaJmKLgk9cm1YnLpe1lXYQebiyaJ
cQPKguzyMkSj2DWg5Rog+ioXIxcAgl1caugKODcrCLw/qnqO8sQI6JarUL2P4i7fTUYfmBAyE0dG
IoFG3288oY/J2J0LF8eGkC08BZKlhiImwP+BaKxHz0UP6zU6oM8izirmqG29rzm4kcUWixDFfWa9
EJ9CpQuG8/LthONgDxMxjJBUqUQgrQyNI7LBssFa3247RxRux6MAb8rdtcG9yt3Smp3D9WZuDD/n
KxTTXP2NYARcLJ0i2ajPK4xHjHhNV+AFBz6BSULb3Z9P65Kf9Dn5tYlUi4Drf1RFSSETbZmiRncc
3R+icUnYUNF2japX1y8Nz3mAaKjT9f4AsLaIu0GEgbos3Ogwzj+hCjoYzdd6Oga6sc72kp8mHTNr
+oCRsMYUwM4Dro520bmDN01he0c9kTS0/Mqj+N6Y6bUEHhkksZHlyK0e9PD+nbkkxIlAfyT72+Ve
8rclxqlnJS8wNiqfVOidKn1ojQ+oeDWJPKGFfgqiW2qLJ3VOzRrcmo9QwKxpG4qjaiOgNh2QfX/H
4/YCCLWTHf73NodsTksY5ol9F66VNnOflJLXMu2EmaTWleR4Tk2CSZSr4u+ff11HTrsNn2QGZiUv
NJ3P+Av1rZIESA1vNq2F4PzqnoXDIGyMCr5Icp+Kz7C3UTbxl1b5HujSJNe9LiGf/DVbBrn6QGyu
QwQUjgzidX7GP/UGga7aqZQoJfbvGS0ltgV6fVW+PU1REjWZoVr3ofzPoKcwf0KuAprAw1B/3uJE
gmmreXt/E98bLKq01YMYLm+Ja9bzMvIEQfgKWyLoTFOP2jcI9U3ASuMqXR1aIa9KJOygcb25BzUQ
MilUbv9yYZGdxgj3VjimYwjIK7ge8Cwu2LTbPi9/xXCHpI5GDX3DLW54tmk6HRUXzGFOYpipi7Un
9JF7/OSz8iQ1R0T+Gf40ud1CkRNacPzxliC4FJS2Cdgjhujp/u07Ij6S/IQTYskn/tKPG6UtLUXE
3HE0LMVwnVE0JfBne8d4R1uy6WEVr9ChH6aK3NESch+d7u6FePrtxmrrboFcLrFcmswCSfuhiga2
OXyQkm/SHRY5x38mAwlKJSa5kTR66pPpW1hsRa3qvZbRT8B2lQEXMITrPoKYrb51UxtkyCKeFK8L
/v3h0Oeizt1ypJqiOW0CHwvG5bHDkyJ388+F2MwXxTOm+K9aKwMQ2wxkfR1A32r7zXi+7rLkoRMB
UUeO2AT/ksCO+Bcar92wsTDyKOjOUvQLOkaVHOofKTnMHgI/Wqlq+YVkCyWdeYUZU8dBJHbQaPpn
11Gi81ciTpCdikt9RdX5R9blZoxTugEXjTTxGLD/dtsKmSd9Mk8ffF/GPHLFh4BX8gs3hdHo7Ap/
17W0z+bvEA7zV4pD/UsjaHaK0RR7n7oKVPLNMDJ8Mr9UjzjaxLJd3LCuYHbexXO+95CYAa3dboUl
T+MpsxLoSW7RbXOl5XU55925OYUAKYGhOgGb6vmoIa8cklmIhm9iA/M28FjdBFgIxGSTbtS0GFUw
zxAm/cEn4j/d1KC/HLi2Q5oRSb8987r3+PAW2VXk3s5xz9LWidw/FdYv/7AdEZxxaB4gDubhhAIz
uVzE0URI/zk18XVmY6E7y+MPBc8UTphbL55nmLJAVGrLn7j2L0TXBuNbMx9rkcf4J2kCopC6/OrG
lnflXRRUP3s1mu2CCxlqzZDp2g+6cLYGBhtXv6yJO9k4QsPHNRSLKVuaMBtI1w5W8Re6W1XajEkU
/WMOx/Sz6x86uk1oYNgzhZjPcPZBbL1zbzeVd/lfOypH4P1qgwe7+fOcx2kDYp0h4ei+mIZX0YeA
gX4CItNAe0d/4DF/oXfKUqbT2GstSe18qmGnaXVJJ6k99RuzgknpUdn/V1VWF+E5Bju2A/lghoTT
MP2iziBJ9lBWWSKagWHja6MdG173CMGxYXuQ6DiUG88jofjk288pcT0d7B9rmJ1cjS7u1sAUU8xu
48lE/vmpBh/DSUSeknzW+ZnlCfe6LNBYGootXQpsEPA0puwWKqSMtKQDR37cohpkZl1S8yd6y9+E
oGULyt5zWjmkDQNcrV7N/ty4gESftwIXv51G/TvldgOSBykV8kC1QjWni6FyygqPZTyYYw1s9d60
pb9zmmlewP6G7HSLMdnpX+CmpCC55NmBgQQsWev0lU5gDEQQqGG515XVOLc6j493K+yE7us0ZvDR
4onHuSBXOdIQLPzrUkChf8Otw/9a+H0WJDksGFi7G7ul3icpM5bS1+CRDtpmnE2g/k0utoxOHtbd
LsKdDqdjwWyQbWTHdihC0wKpTykxFvvBnPBDu8p9R/egvIS35Cj6kjLH6N7XgKUWGmj1VvscCt95
34njH6zywwKyNWjLdcr4Vn285e3Bxp/Xy7f2tZLmuQp3oqRkyQn+SKc5rZFaGYW5rXkvuGMEnZsD
BkkYo+Gm/QuaJtNiQCLdS+O9ab8VP7ZSYdzwzMwFVU8aNOVGOzVw69mJ6NpL+9HoLkp5QD8xiIP4
KOQ+8IRSTXgfYhLXzWEBquI8do+iC/X/bB1rTl8S83T2Db4JkODTRynGXizOVet4a+3e7p0+nXW0
J6k5obvl94rEUfsbESdswgfQFFaXrkTDUadnd2ULQjldUxQyDSli4Z5Mzr1sIZEc8v959YdazkYa
ebQ5GkqlUbdv4PMWA30V9BaPbLCUbFwW9xIaNt7aT6qHBCwmVyMWdTlt3yIqTuP9sBx/g8f9TGQs
aHdIDgtPn9VDC5yWBByM1TkC4npKnRzY/X9brlD3fU9lPZToHPOn21NtSX0hxQL9CbDt8Jne0Ugg
qsyhGOh7x1iKANrS5YF2RsjBJjvFCbVI1lVGqkSvfwaXSpHX3FB4RJFVdMz60pcIxB9GODRAyl9y
lGmjJZZrzYGI+1bViRHkVGnv5fs3mlaLhRYkd3oA4Ua/KToHJXpXj2xMOCgCPX3oSJuyjyHM3GOK
jlCla+6ZmD2tV3dc3mUCQjZzg1UAvCo81gXZsWu5LPVDWXm74nZymABNQpWCPDGbddzz4oKb/1wS
PrO9Ckli1eLQ7Rbholklnaqt592+WkTZiy/CL6ZiKb7m5mOxtaeu54W8V5ne8Fuj7tS4zxgBqzLY
KYIc/IAdfLdIR5VdLPShF+ziKI68pC58c1E1ZsH+BqtK0Vp5tVKY07XrH195IwRledItsHPWv5P+
GxfjQBBoEIG+yqHaS3m3ImLBTZ4tJ4cWxPi8h62WFbe3LFHF755+GpTpRCzVHkHum6/+rIyH1nQ+
dE7+3EeoI+V5BhvVvn5dNcNJhCfWOLXm8lu1MBx4xUr97ZXB0ezcnH2zFConpZrHbSjX5k99wDXK
EJjw2NZJHynLk/JRmGq651W4f2BTsoT36QKa2+AO2ADa3sacjtM2exQzHCDG6RVfL/R7qKaSau8c
FL3JvYfTJO32b1CgoivlNJ+U1ELjnUTsuhhLwk6HGsP33Rgwz0pqBGFC0JkVq6HtNDkN6Ru663CG
mWWq7ckbrEMHmooQd8vNIgd/6rS/6j8VtEJkY8eqA5WilyBXqm3J+xpzTtnLjoCo5MLSxE963M4O
pHFswjkxIfdoS2P8F39dlFbQdP4bTYI+L6dNLJtbeexj7zqwYcKx+0YRU/XtsMkY81/Q2KvttSG7
E3QHaAbskGwMbauCTAhRfpAaFzCNoj3rRQ8KeLMXVk/uUlfHui/KvE32ArVvdufRfGt+FEnJCs0g
kYyDoC2AXOZG9kdtVGKakSle92NkJO4rU7OstuejxjdsRKuTz2wrcJiJJg3TPCd/eB7VqOgHOrS4
yK14Xf2JgGoDuOUHV/eayfpq4XJfkw4vo6pVF96soPW0NpG80I4pk8NpO3S1khY+/zWwi/JKPAE5
ui0Hm8ISCyxG0SUPPLapL9kii70MQ1Vnuqg6eoMXQtQ12gUOr0fhyVFZtVokK7sR+xGQQrnvZvCt
1ztE52UaiWRlju7U2D7Fm0y2TY7obaRXOs8jYGfiM5bO/wrxzRppnHnnLG/5y5ZB1K4jrO3R8rbY
LXtNPLUCy1Jcv3KYneagg+4bWk9T0/2Z+j9EU/I3ixnropxlF5BIN30fsebIJAnqw7XQeXOfhNJo
FrIuqtFEvP/LuIpmmdD0v2VBc4C8M+zSwRG8mQaJJ4CyERxt4jlpPOSwpmLuX9UBBclTH4UDCITc
Ybxx2GCELcZDFF/0vY0jhDFCmgoXt5Ch5ss0EQAWkpN+nTVeDtXfFZRRjExTEbfbJdDKF+jN/C0C
sukFp/8UgPpP7jkSS54nEMRF7KTFQn1rGFEtUZHWsIVbz2W+MGiCHSB8U73f0EP2KSdLFF1iD/OJ
xpev+h/sNBzRpa39nMIordprKldHc8O5sF28nk0qPuE5YlybGfSv+efFG0R+MRwVRTvJSS7PcZ4C
hFZ3mt0mVtdNtgS+rF0jtrd76FJpYNtJIX+yrr36cTON3BzW739IYw0C9WN5FhFnjR+y/f4PYDA0
dK+uXidMZaGd/SXnwuuLX9E+OA1efaME62y8v5gEaG5HJ8ovjJwO0PzG4qzKL2/3OmQSm0M2Y+6/
g2fkcNBBNmtb3/cCcGpeHWphgfMmK03eJ58QxZN4/mq4upaTuVFLZC7m1npGibXKEnqTZonRTPrH
e7iFLaJCTdDnjD09hxD0c7SxQxMV2ExGWXNJ4YLPtaOUr+GLxBabbUA5/JhHOI5ffkD6hbC5e8y4
kuujySu2CIz4lYOnkhnin+G/ew9wJ6zR3Tx4CkIVXh3wH/QfJWo+jPeMg9K1hBUpFv2ddmvOpIEE
VTesAvJUE3USwjatydgbBnvgf6v41fwJyQAoF01RXf54LpghSK6V4T18q+HvY+XaoHVZS7nofy2E
n1MHzt8xFU4uVErlZEQFbSZy51+LABN9FvD3RKsrqttOor3bLBwu4yBjX2wToqEDBeG3M5F6HGSS
ZvcrkyeHrnkShwMv+YX0cpeHNgOrOepnL7zjGOYOb6ojSYKTG2vSGjSiRZqSJs5nlJm94zHVvXDP
erOjZfM4Ws3lm+Q/Duy5SUiWfpr47Rg85aXGH8aeYwndpc3pKRpHLm17HcqGluDAwjk91kCfDVgX
AIuyf3P574hGGnnlCeXfTPKRYI0nbD4ueWhWXkeCx5qP1kSF/PFcPCkOq/2G4CWMmUGPnCK3D4H7
B0ifRl9QzgqzP8PhefIi8uXz3Xc6Rhj8ClI0eve1OhdisfclGExkyH96rYo4SfBlVWcYyv2aXNcJ
mF5Fr4xjkoSW1b8uF9pNTRWEzZxkfc40IhI17pLwhd8rLJWwnGadgIf1aVzMWiTQIMXOf5fO15YI
LWGj6PCTsxjFGhDRq5EqGtHWZZ8tP1FJMBHorY51riFlV6vt2RGutq3+I5gNMnbjTHlT0F4j2Qp3
Mc94PBgRX+xCqycjnshhPaItwPAsEiPOQ5/qdhEmeFCsHto0xClhKUE0GJJcvX5A7qxPwTTjk1uY
QVEpNDY17C5FqD3snyd3GefZh18FOCbY247IpPdsePW80/eHVqnLhRZoQ8HCZ/PiPKp0hd/wyT/s
K0df8lbNkYSXtkR+ksuiix7sjilc4oxBNM9eyQKmvxRnpwTBMaVzu0VG+rCCclJ0yLP70dklPVbT
/K9uVVlE5fMXHKJo0AqTcApB6gP+MPZLYbw86uNrcAFlr49LeZReIQKUa8xU+iai0eAR//5tf8Q9
ok7VxDBlCMhLr1AHbIK1Qh5IpOADy73lGD/CQbEfbr0PEaiyzpyG2IVk/6O4q3AVXN2mlbHcKqhW
r2HUsZYb0HubZiwHvrh63ccmIImotP0B+ir7B2xIlQIW5Nw1y6ysVSDaDH8r5gio3MN6vem2aXjJ
kB5+4iE9DPZB/bOGTEXTLG234iG2zvqmH6QqT7xT5U/zHj8U8/vUICwqmj6Y05ptpzU/96PRqd2V
pl+VZzDbZfUmojj33lR4uT6QL+X6q1q7FLeWugz0wHaV3PQCvHiKWcUbDVQbXREJ5PsPQt8BSHHf
hQwgEVVkbn61NSpUvEm/DTs8bRQmwAefaHMEwwN7qIPkjCjpUCzQZirqbcpUvpc0Ak3JO3vsIlH1
7h5llUtMqqiq00OuLoxeTFzsoaZaRD7kivTVQEbqHo6QuhK+x+sNOhhbnTbZ5YpbhtZudA5M/Q5g
4WH3Q+MRK+SUSMMn+H7KIPo4TbnqBLz12ycxFwmOuRj+oRr2QGiXzhemXq4NxVSrqRF1oifsiO+w
n9DyldozSN6703ImbDI+bvESlLSGSiejqTsSYUfJys6DiKGbSBcrLPcGN1tnIWYaT+Nt3yne7VeM
VxjKtFiBRWpM9YpOhFbOE2aaKY11YGM+nHu7nvSzDkl7xDqKe5kqaaibz4fyqjvl0Ox+uCum3cL+
VeWiYCI4Z0DSvaul48grbsebjTrT9unQUtsPKnuQonXuuLMo+xAVy5gfnhfXQqDzpzERdQNhGgll
hDgTUUT1byQAli4OYkHvBtJUObVPVg3TU2xnQazkeJ1oPM5hi3AzTEbsTNd9XNuUobo2vCd+0K87
GFdd4kR8xS0pko0qOlb5lsYUAFL6K1PB/mGQZMmfnQ0JaOuWNPs3LSVKShDivAvWRja+MB+P4SOO
UO9UR4tqGMd2h5iKtlY+n06YxIDe9eMiinMnF60kMQW0AMGJa190S8fPnYjLjyj7dZ5+dsR6cgBu
mBdyUbE7OhIG5bQnvHCxZ1BFmdAW9xq3tOvCeo/DqcHrprt01fIzY6asKhtEYlVmlGR0hT5ITXE5
uUH8DEsPdzxCz3rPa8+d3MuJMG6QEyS+KbfF2a/bYL+QtVXzEqWMn4gZLeQlAAkZYwUmmutl6WK/
D2Pvmy6QtyfYXSrtgBSSj6WRwc7UaWtGVzVKM9hUF5vomVRJcPWnenC+PKHXj3QNztD6x+K4gd7F
p9NFWL7v32BfH/7OCEJUKQTZ4mgi8n49irG3wcqliiRdKSfbsiu6jVnYCDtDF0/fZG0nSXo4rNjb
cFGP30c3+v2E5ZTL5+ahF8lvqiIbGYZEnjchl4BXmz5QPJbEWswMCk75ZPPDFPMqNTiWbOrzkhr6
6DX4egrmX/45VJ1CLdylGtivR6vhiRSoRXKJG+Sot25fFn5uqLS/iJzunCBel5CaM+8FiaHJDYEz
vS2iXd9zMvLNNacjvYXT0U+/SvRgl8+4Looov+SxemkA6+PIwq7pUvFP5v2qdnkqQH75EYWN2/Fx
JKE2WhUGNY6OFkHNZfps6AQSoUjaIe2hK3j6fWlaRYgyLjIbV1+GvW3ry5aca0s1503dV26X7fXa
2PUsazcOvC7gstrz7oIXpE4ED0gFJmeZMB1GcT4D/yNYYMtprsFBfQKkHKUgOI03C6roD597QEdH
R5Xc7LxRfsLvm16MlTWoY0AeL9FJG3glFBFVC9olKl5IcWg1Q3Wijk3p86sJobKX/4sKXKNBaTL8
ZWstb/bXHvX5u8opI9bu68lC4vyikog7a+e5gjCF9xQEy0zNvYK5RtGuV5R873UK9EbFR5Reuzrp
gk+meTMJR8C0lcPWLVgGw+IIGITzzhW7+ptM+SlqkspYCljTZy1raVIsjlEjODaxlr5dpQZOVD2y
qgTk2GLR/0SZD9NqtTAwDgIA6OuQ4JEHeHzmrKX3k/NCkKSxmcAlFCMkuFuDZIXtkdE32KS7BQll
3TG/JCf8msBnMktxtif56gkkpu5x9KmKMnDD/rzVNvRPQNIiaVBwXS4QpsycJGDE+K2elzB7ilNf
RTdixCUNlD60LkTBmCRIeQxbX548L1v81VudbTeuuQ8+CPjtIxURSIQEGymcaoyogEqLPjKSH6zh
zgDVELVnbNBPpFZr/MiKH0DuOTfJDDfxIqqGxJilKaebZBg69vo2qhjujsicfEwHv6B1yN5lkIkt
KGsS6i3CUYbpEQzfdZ9KI7JGlKwfM1jQ9NlKdAQ/KC4UnEKbz46MTCxrH4xqG3ZQS2CaA2gkw45U
1G77TpNdIRmiBsttp6dGx5cqVGrXvCe4SoJH1ipUiWj46bjP5IMabeh5AThM1iFKKIVdFPMNEsbR
fApYG27Ys3TD3H7OJnprb19oKZBYdbIH+PkIlGqNG+6SD6V05cZHan/lGdZRCk1OEphovUedHnKK
VqQIbBPROglSWGm8EeRs0r1NzBUfTHhLait6fWfwqIZ/J8N5xtOj0DlbSpWkc3k17Pb5xJ+VvGWm
zITHZTtNPks7S/7HxN45Xajbw57A322kh6m+i4pm1hUnfQf+wgPXCXrCElp7aIz/mmbuCDzXKI5A
xj6CO73CP4q3MHwaAS9sVjIK+e5e99mu9Jr8LJFDi9ms+6Mhle0W1MXRVnmJ+fvPnRRK2mymhjDx
jRc7GNBpbmz1nBHmAVL4B/b0F9mp9tWZpDD9u7I2UkHBw0WfGsithYsmlZ9RZ8a6ZmO0iRDv8k2M
GHq2Aj93O2T56zYxPVVD3P7ySBhyC/VTNKS+qJUQ0JbPBVS4+hHfGJvVOAmHBJxOqkOLV9ke/Q0D
9OUAsYmgmBqGIbZYkjLqk0trJ5IOzwA++0tyvPknJ+2WoWJRFHSe3nr1ZfqlCVnIGOkBMa5w3oSt
c9I7CGXIQQEWp9P5TZI87pX/TyuFxqufVxe9gBGb8vppBDQ/1tuMeQHVAH1Vr7XZSXJEJdJkYzRP
vnYg8oc75FIap00XduuLQMMLjlk28fIJvs0x0qByOXLbyWvwpOhedaldKH8v3hKRAdTjZ5wU4arr
6wEGoQgVv4RnXLpDr2F8mRvZ6JTu5+X4Ud2zPVekuS1DqV4XVpG/FuzF7GwQy11fBWDU2sNuQS31
LXokDkp+FSxP7DLrw53lA+I32+hb4X6P0GNCuSQ0YLq+g7CflXqH96yhlwyL+TRZEqiN6EQGr0kO
E3n83PgJIgVLqaN8+mkjQ5s/Vq1DApUscChxWuak2FZBj9oAxT0UBnyrUdMnLf9h/6mJZt+4AQGC
6ez/tFj9PuIARgJ2hesW7q1j19PhWNDKp2kh0pGOEFUD8gaplNbOdAWIUv4OavONgn9yf0Z8yF0O
UEk9LM1XEWqMVcx0vg7kHFXBHY/Jm0BzQxcVU8qW/CFGTefEmQwE0YilcSlLzoxYvZsibdnl/ETS
PmS3bSDbQ6uglFsIjDtEXJer+kEK6Iat8E0jBE3c3OPLV3v/sSbqMtYqiPufk7oxubwgUrozk7KV
9VEW1GG361WYGRFuLTl2cK9trdMN58Cw7Zx9h4Kqm6ZY2mK3lJmjgdMqsmUDzZA6AtMsZBeYoD/b
uAAdEob9r90FsG8pQrJOhasbhGs12xJPeKJVDXUYX4eZ+RFh+5BLssrPTaG9LLXIwTYe/CK1B0Zo
1vOj+Xv5zp1dtzPzkOFUj4OCqnwuKy6wdS+bRKUJfps2WGlsfkn6Bt7VFfZq44S/NfD7tQHxjLHo
XUKGBK4x7xACOWey5fFf3o2Ncn1hSOg8HXsamLx7U5vsY9dbwEX87W0nIM4p7EDo11/r7YQLEO7Y
ridJt92wPIFyVClPcNE2FWjbcwifsNAZrVbKkXEg2aak9XvkKo1S5i0Pi8UljyQScsNwbvrAfqzj
oDqccEWnxAgQfAaBpEfGLhT2KNzCqqh7N5cPnQwzyUGuT/E7jSdUl0UVJqn5Yk7GGzFMTCyUG0Ku
UpnaJrB6iwF1Q98+qTNQLl5dYM4o3n7NCvSlNASZ/jLg98fqZqUL9MN1DtZrVjZifzvvIVTY7tzZ
WKH33vTCfJlze2rgHiMRE/Fi+rh8hIbEiLBB0vokjcmjZdTl3povWOqPetXvOF0N9+IiM38X51gz
oYI1ccfd/HylQsogrQD81Ey8JerGrCb41D88JXjun/d3+NH19RmbslGRowCLkAKf+k8IlRQRmSie
ZAV7/TgsKkWKCN/LJ/8C6qIj0Ok/sr5gJ7whWmYfCwDGdSj2bHoWXRd3S/cJeXhVD1fIZLsMb4Xw
3DvbNQtXRN+VEd1N1dIv7KDoRxCS4l7vk4AEC5UQTaX6yrRjd9CaCwubV5w+KIgjTsg+R1Cq9j7V
F8PEXR8IKwzkbxYpe22DUe9rqKWBa67fjrwY/ltpN2b/cmOgiQGxEht5bjbw+HAHGWAqokg3+JZ7
vraM2r8Hkkx+GxdTHe9dAsWmiIclEelZibONh5cOZ+1+8FJJEoBB/H9ZEjYZXrpUC53P5tyWI0KG
zUWB9U6BIqZvy7z5AeqAjWjM4x31kIrXNzAKWCJTshTpjPWc5Yh5cAltuBO3AQpBG75tKXkRIoht
m5mdXB1lK6YYUfaK3y/nk66sMIen84W56k+s3YkMT1fY8CHyrqFaT51P7f1xmirQ0bAZZo67J1lx
Vb9SVSvtF8GRcg/0pyInRtqDCxZyGl5GmqgOyMONq5WkiASKNqbSYs3aDBqL3+rEUMC5BNwmZrxJ
q/isD1S4JPXF9vQTr5orKRMyOfd9qxmHMYuBl5ge+ZVnWoihEolEC4IzAK/K6W864LabGCyCSm8E
oo/fV1B4g3D2IZK6sIGed6E+/8/nskl3s+V+61Drk6+2uGdjwRoXE6be9Dr7kSbjQmTa8uXmad6x
OmssQon39ujEg4qTyd9ISl1TqSVDtV5Mk1ODf/kSbivbG8i1xauEkxFHQaQVwDF/qGjrVCpBHAyj
MMaqJszQ/aGDQMc/SsmzLUYCSm1Thcj10vBVU2Sd/SwE8PUYc98WhMQZLJCGIzUiyW/cBSl/qaYm
KBsX517Rp7KKJCryrkEGMUR5uD1SbZvloLuCHgrqPTfKsCIoBOmPP2ZIOg1WntXomqbMrJTperrN
+nQl7hp2MFqXiaw4Y9XgybuP3e6PeNhwNc9uiWNdNiI3NkYvMvnmlpkkAfD6385y7n0+0YQ6gKgQ
pdFh01MbviJoXl5AH4DjniI4zqnkv/c8BqnI4Oz6TgZuYTmJulqMqtyH/+nHq1agTrP4SaC9Wr1z
fX+s/l3a5fmrTRplRDydQbRISNvRYO90NUyLJKKU0FnjJIIenXl/9QkLcuzdjQFD19NDOtJZbw8O
Oyqp1DJHcdkj7mNwa0FIpe9mMz/NXF/AmQjbBEXJ8WdtJapJxUGnatuMKvH6/xseR15mltnTGlqb
KGpT5WTCq2ivjpl7LCN9lCGjh3u5s95SzNrdQQsTg3H2H4UzSLCT24C+i9IWeElW4AgGiWECrcPW
3Qco/nx1PbboORF7qcS4EYQty2NjcCk5KDWDcECgya4p+OEwo3TR0uJVmYZBvZxCjv1StqqRd7WZ
1gLiYOEaAjZpgJu6c7sI4sfSTO86enmwDgM8ZfJNKH6EkRyzw641hQYU3QFWERNT4kq1vJ8M8ndH
EYxmn/iVT181IFI/X5gBx1AimYN/r6sgDe3lbk8p8nAdmdTUwRxgi1HDA7VlqAtSNd0uFmOyfCeQ
R8CFaOXdk9VNSirGJPN8n5VUvRuW4RoIU8xBNjxAT+Lf2mwaIbdQAt1XrDtB+Er0U9nK9s51UdoI
VksJSl9e61l7VjB/B2M5+TclABEePB5dY9SvFREfadApBVMr5zS7INBsXfJ7We0wsqHfLZtQJ6Vc
aDwBXSxEqMqs/5+WOO+lZJSpxiGdHjm6JI8vDjsHEe1qazuyvhkzSzX+GPSz64iUk8suSAN1xBL5
evAHG7i0JePW36OYFHgj2sSWZ542QB0EiDm4jNK8Cg5KDKptSeQ2EpdyxGUE9XBdX6z/f1HPtK1t
IqYk4PGJNZm/7OCb9THibxT2ebfdQObhJpK1pkB5bDvlEYmnOCQWa9GeNKbqSDqsqTKKsSK5H0ZT
/ZJpWe0KUh+WxEDItBg8ZCDChKRlrT9WzdcaLvaFUXMNi5exC13KS4fFftvLFoiUXyMf4wQmpkAz
PwIYsu5Pk+CSAYVA1XEUDc4WBgD9A3+N8bsN8/OhoV6kQWsY/vNPwEG+uaiWFfyev00eJeZwm1WH
V+e33XuuMjw2eJsFXbjggp7b/bDnqnnHKnuwf9SX26aBXwM6Gh4hwZKnT0AbsypCn4ftbMA0l+3o
NNOj9HDMMfpN52atgGGEbnpZahr3yNbmvoxeyMsLIRhlAfJBwVF/c7rEwa6s3+1xOsHlyIoqC22Q
00yhOU3u1w6r7saoGnH0BK3tuu3OQtWUwYLUsmF99I5RgbttBCf+Hi9+u6qbuQCuzNF6HIFW1Zii
xHImtIOVhitMhqSrDQmNWYshVyVz4PMYVJoL9PwGOoBPKLW56ArCoA42jxmWIhL5suiDldNpGV4H
MgdoJxp85Te44VXYn9xyKLx+5QJVeNJI02a4NU9JRxYq5lWSRB2j1/93A8Ukjnnp1xfVK/9RzKMH
63EGJPgsIWeEwmonhLgwLRN/HKxkBS25HwfQAuAU3X3b0A1iNcswx4Slk1H8caNuDhQVyBUxKKuc
FVUcaB8uzH/i430b914RSq85oo/wcHMGB21hqvC7ioMjBnxk3P4PsSwLZ2Ub4AHfjTckXw8qXDJL
P4fOyjf45HDa4/GN6X3i40m4C/Y1E1/VzJ6Hol8kVdOW0F4I2AoWFmu9HocmadOZYzj6+d1vVcGV
2Ggdt7ou9uYd8dEaQeuOuvGQx/YOBqjrATw14iTRVauqIl+NFitHpE7ub5FqTJXSR2pQW/kwkWkj
eixmFJSiEWG3XDE6Kw8o3+tjaM5MYJ4KzifPE61TxYzQi5xGgDVhQcelQtovISBXHif6KxQzOwL3
d3bHzUvh1wYuLau1b+T4mapECuy46hH6IkfULu54hU5feyhX/+WoleuU3dAcobkIOWiQnXhvlXbS
2h8T/pZEKuUOcB1Q4Wfu3raVZBWld3QhzMHStJgIzSUoYbjgPiKdm65YYvv7IzmtmNtvT4QEZwGG
N4s4hHnYXwtIAdSvTjgUR+6fEhVFwkUkUgfHEwsmfVoS+5sFOQMxKYtllwbabbZlA/5mnUzF6GXr
jnLW7PYDS0gKwgybVNcADyoPhNeedwDYk+QoIlU8YY9rxMRlndzz7GLVbnpaSe/c2jITCWd7zNvH
glk30gEvq+zSQr05LidcDHfJmkpI3RZLc9TFitTw+2wf6qI4bNxp38+GAyYZH2Bf+waYp8a4hFl1
dcR/8K549uNSB/Eq1679quVAv8i8jH/twwUkotnahw6jW4M8gZSDNeuRBFX9XIHLVno6nz9hsRt5
+6pzI8e3un+vuz+9RxQnsFx1SmbFXAf2NOf5WHvtXxJrZO461+7nIO95FkUBOU7cit5TpzfZQxvA
3N6LdEBi5ptZHOFBdQmPldSTbms0sq7l5j6L/YpUmtEDcXIMTVEyk+TutMF5Dutl+ybOuK6QUE/3
0/HTwU+jqBhzlLUFgEFSc1I6uztaEhUsK4hCUIpiXnzC1Eoo/0M5EW+v/LDfGM9eFfmumavK8/9Q
BEtuuhtsZOKI7pmmeUQfk4qGP542f42XZXYiZq6L7o5QUgI1b8OqROwpwa1FBVo62cCa9LSnTaau
3ShY8b9EpZmmnvtfUGp1eMjIOrmg8TpxTHnxb5BIIOonRbobp+FJZajldESMlquUDqiOBdvOcPaA
7UkS6WNz7ovlg7eA4qf62czxK8hA1Ah7rcqRM3kpO505TeZ3to+t8NteERaPWeiGdQfz+CbjzuF7
qXiOq3D6BA+w3/zcxFVPA1cOhE3xud9lCucDba3dy3QwB192Aq9JEeUwOd6wC7YApuMV9f8wqLP1
fpsLKtyqOlpTqCAG8IPQTbbWYCJ5INUPdfC2TXkl3LGkEZ0ICWZcC0gsIWrZZdwfGfBzPkhERa2g
2MbEiCj+u0QiuN2ZostHxl2kR1RzEWggWrEK7zrqheS2S0GP2xOCt5jHPN6/t9CvOzKxTj1OGfmO
Jwg8ZVnSwIVDJwsRNDFa11iob+8zqS+fkCbHLOxxWzsKYlHOYj0+KpaltK8PiGtGIedcsL4sFOvu
8NeMfInKy2WSTEorNpWpZBXGI0UUINLe5dDD3RVZbo3Y07yl/3a35EK7JAygkHBQ4jmzEE/P8TUH
aFNkDzzYdj6re8/azUhh/bofexv0CGg9OWUMB8ZemRfKd7sF7CbdpwddMaeAKheTKbx8AeiG6r9h
xow2mW4rtmWdfTiBIvSRizCZJVRUB/BwWu7WfFlgqsP2fQf5kgxEWy7TuqFpn9PeDA00fUBRqXUE
w3Q1TI5onAstRShu+i8MqrBwz38NZ9jzdQCqPmg4kSoDTvKcG00b4C6POVDL5CO0Efr4Ib0UrV4g
JwsRT0uiInCMkT4LC900xvCTu+seqgxGghB5ncSIfxkpLO0BMnYY/3yz3hRcuBUiBqiLd0KQaDqf
z3PLB3/6c2C4cmV8P3wzOQmJibvu52scBy5xfY2KRoUECOdZ0sZoZiSpw941GWz0FjRD91T83iYJ
ckwEad4n5lvsEwFdPNGf8LSmCs6UOVYGkIZfdvEjh+B+TkubSTmorVllnSUbdZsZBjURaRAM/Zy7
z9lkKsmwamMlVwbd5XmJu8mxgGQwC/ydJ32J2OXHS+uJ1oEpMAAExHB7eMrDiXhSEJ3sJdIUs33m
Bcd8bJFgRG05BT609YehAnIxbbp9wPW0wxubb1FHO8sMehojh/aShlVx8hpCN942Pg9vcCSQle4R
0Ii/uwaNwNNa3DFOgAqJv0qV00h82g1utPUfk25zeztttqaormMWcN9OHvqyvr1C/IYvoTO/uWy9
Rez/xCWlFs909r9MfqdCB491IEXvLAKUWgy8GsOKfGpIEuZT3CNRQCcs7BCpkiPoEyaASIQKRZUQ
z6Gz0h8Hhc+Ud0Glkrrl2LPO1tBHtiPsuHVOC3ncbUGFoYdW9OTK4cFYg7OoDOBZw59meozykd+q
7GwrlMkCYbOHOyB3QELAib6iXBbn3q5UDV5Zkj1aIB7bkgwCZpIG2mLGljJA5tfsA7YajWYXsaEK
Y7gwAZ+hltgpEJl70GGy7rAt7S3LWQm3JSVBPLouCuh3z9SefSYs0JBTYlML0zIbrVo7HaR/5zRu
HI/DQ/3cb1BX+XTKhCUi4FQpNDH1E7voK8m+DdzMoEVzw0s63bEiteC2MgMtzg9BbRcG50y8E00k
lbuxjj9YKlreGV8Cy18r//Z/3dg7QsXTP7EsGNrZcpyK0oJjNm2G2EPcAijUx5SqMbUhvw0u/SVY
z4e8+lQaKGKQgqJz+3tImXgwpJZkbN1nqvcwMfQnfQkFrgtRIpsyLHI2SDagJ0BhlKEokY+KFwT6
cIW43eL8qmadUXlodFfPM2UXOJF3ev6RYItmR+V2bw9YUhuNkxhFQse9fW7ZOQcH9KCGvt9qSBWs
wqmAIzGnavL+2EHBYKROSoEcn0ORDkRTWMi0U317GIi0ArezNorpWwSbfV75q/v4VfSZtUySuhJM
VDgriDYmQxkLdDWsUxxKrQn26lkX8noH0fk5aYZCRlTEtZP3dY4/TTPFdYQImFaZxanmOhUNjm+0
ndlmEzHzFOjYgPXdl8DfSu1Z15M7kFagn29JHOREpbXFXN1x7tRwMOibxMrcXEf1CYfYVMLn9Maw
Jx7qPOlom+btqXiZBaPll2sjyTBbb0blaGE6ERzLT0jKLqN1PHVtKpubbOMgA3tHsOu9qFMtFSsL
GH28W8WqJd/WtTpA+q/2V7Ie+IEelt5ME1VT/LntS7BqepYyh7J4u98Nv2AVhv/fOYXwyE6Dy3eF
7O48ERgjLXREvFmjfqIR3GZhhZA7DxUioFgSI04Zo5VIGw+SsDDeUIumKpmxbLr9EeG+VYPZvLC3
uPkwBRTTFJNqaF2wk1xualaJ5hSTPiiJ6UlFLZYmD/aPYmDiS3mY38ZN1l6Oi8aGwUOh7xMMRBvx
Pv1n+LCq39dD6gyJZxS2lc746fCYh1MrfmnYtYQcyQYku/876FkCcFxXEf7m1vwwHRkH6nAfAx/4
/hQLHlYU5FruEAX6IlDtcegZ1qwiNyCkemw9INMQ3uCZA51dFUdDNCNzhUtJHZzZNrnaDoKFBnSA
PEVFOMO3v8d8zn6wBJ3ZidtnGMGZLuKAYvxR02aW/AevgcnZDwzwBd+o/ACOIwn8SFzU6WRj/YKI
JB5MY89u1X0aebNAxiwDIpfSMWgIi3f6lHYoK+eVQnPILDY/EtHHOfx8dLkIXfjL7KynQFPwbpsC
aiyszR9tmtVZqw7hWxqxtMltAShauYeTYlbKiy7WxeypMW/koQW7rAnrObt5tdd8VSTgTUhbB+Mp
fft4bRDrgQaQNG8XRHYsTeG0cV1DaQq4JI34qe69OcgSsWy8Cf0y/YT1eh8l4j82tPqYjbiRJVT9
83uL4JdXcNYoC7tOplX0go7m+B4RKRbCLHMVOGNix96ALJu4rOwPgs/ybOt1Q+sTuk7JFKlKeilq
x1lwLpncDtW9TjuDmsWzv4eBu3UsVZsX6TYJYPrlWVk7uLfR+ucAeOVkIzmkZp/FLsyYEb9j3Vy5
Z/5TrbwxgmwSfirG9pjQniQ9nYfqnz/22zdiWTYrAiwKhHu6rUPpyVVhiWeXBkZK2uFPCmQxEz2A
xrQ8l0Olz8AHYpjMLUGFEcu1hjR//9huLb3zSbjJgxBUeWEK0rgbOz9Z63is7OnYroXz/SmJOAJc
FmKJbV402sjLfDMm2yCht3QxVReJB0Y300kF4/tGdiK8DvXEAdc+ZZAvS0bu4L8ymKKN5QW2dye2
vPqci3IBKNcCl7n+/mdI4JEES8FeVoye3TRaElT6qWul7Dt19kPzq2ZBJ6wvA4ZT4EvJLa27Pfpm
PeQKE7hLD5gbFWMQvAXopLTuP7NIx5fS0Pml+ycrrMYh0Zb0oa+1f4QGvD6LLZ7VcfY1QcrTZg93
3Q/PnZkgxCh8IRvKp6ktKhQ/GFCgj7LVS0I7RZY6Swu2NbgSMVpFUOaWa43RW++lA181tpoy2pGz
kER3/7GZ7st71Gkh+jUTIJXZ+KAgbGJlFImkPzFy5y7NQVbQfucc8Lg0jNLrcxxRtcb5ie1U8FrK
vfwVXN/FF6uf84D38nBwndRQx3WN9/UA7Ps3GN6+mtPjGEIEqVFga9bcyCogv6WgEBy7TUJiT1tP
m0wDIH12j9Dpygndu4wUBkgo4gAMS2LiLQyK4TX8jsPDU03iTzbTmVC8hKFGNqmksgxF1OcruQkZ
6WJycl/mhWJ1ifGyqalnChwoA/LFMkCF/uugu1eUeOP8nf0qwkbrI3rmOZHI4UWzE7g6e+riwcPP
KDOBu+kmsTNwwvjKzClChLyuWnW5HFZOD8D4o3G+1jcsmiPgCFnCSKBMCpmU7zXyjnm/1VDtYXIf
YRGPkskVBBMUG3YyzD/ZevJGNbGSW4YyuRxaDQXetK1bvbU4I6r5IERThE4eHxwmFITzq744T7l2
t5TQ1zjP1T6EI4qFgGH+JeG666IVb0hUzEscqj99OlMB+vniy2LXrupU3N1Kzt5bk0Qgn0rBJTaJ
reC4WAbO0/tHZ/j64wkJB6XfC656AZWQLoTwZanxEFFz0JORx4gEmS0l5HekutboXz6rRk5sN4kS
IsPMkmsA2pc2ySzohcCCCLyQX5UG1RctX4FgRDtzFNhEsiHZJQuKK46Z+cYQNocpI9mhArrd1B0m
Y9ehq/hguwBK2IILNA+0cMzA3en0pQe2v3gfnHtKoLN2fGw1NTvreBH6f8e4Ueg/fZg4qD/oWz6W
8oZkT1UOB47gNFxQ/l2laZZ5Hq10uPYcnL6ZIL2Abd2KHL8YdFbNsyhFjUKQDsfnIWFvnjjYKJ+6
4v7+aIfY5lzEBYI4/A0+945db6OMi6TlQXBA5ukuabox3UmJN1j/7P+p8DxHqR9ill+Op43PFaII
vtCK5EYWO/ghqSd65yQCTyvbFP9dY3dkPR4GCDrUxDVa3e0CzeKD5IS3vqvIDJSuDJvmcdxKlixq
4mHY/5Qjw0/JC86Cvmk+cxrcMHGFJaenYbHtwfTqDEfEdaw8v4HO+vL8ZQ6h3CTNx+m84Oj/Mq2S
WaxqKrLd4o0aCRG2WhOXi45n4a/4zTETmKA/nl5qRAfZfhgvdoAGVeuTcLqeIpoPDcaKIMDL3ZSW
GvGYHXGnOKbhu99XAU2KPExNz56lquVJb/Vk9TSqH2hGe7qWj3v52AceIDQZY5RFIZLSZ0UIs4SN
cyUtoUZZ0mWxp2w/QX+GIBi5knuN3Y+tjc4ikZl/DrPZDUtHYnSggLD2R8GWgnvZ8LKnuVZQS4dy
DDsKfPC5Dyz5bkb0+QLEiAhN339+23qyVCwO6PwNTXTLvzAJiq4JUDczQ/zu7PYhU56obwr2YPT/
GPyi5kVmSF998ElTLRBq5UaVVAuB+KjlKUYsVBcv6JEcJOSIFQ/ON6ztbveITzumeCE6tUWQByYz
uWNUsDOYhgaHY/X9a9g+HbSav+E0s2cNSC1n+k3GkxQuFJ0khlFCmI1RW9o9ZM7F7JYFwLWfxOK0
rpr3UlW3XT8RB2MOk0ixRwVb+TzaKEoItiqdsRfc4A3MqPkQfcDWxW1JChdwYxvflh/apRpPoDkR
TXYfLyzHWhJ63BmgVa1MYhmIknEZIqQPCOrfud92HE2cVbO84Og1Y9GIb/PIeZYTzg7g5BTiPgrb
0r4kLSfMQxw08oYb8InZv8jLXCsVifZbVfrW7BgYodJsezTGeJ8NaahlgXyfLMnRRAuHLJwA64H8
VC10aQ7MvqdixOWAvS6E8Nj5iNthxL+T8WNbIyJTZI5Tfgy7CqflhdgTrrhVm0PbJj73AvgJCVhs
xJGaRGbiqGjWUGfzGyZt1cxdWu06qHzfpZqEazebyE/6vVEl6N37xDnhP0zCRCAOBafbSlvMaaYp
+G2YNTvKGkWM12/Ael8bXHDrCCU7WAEUFAjsUd/rDFWcrTjFA9ONsgpk9Keu5acFqV73N0YxQq3d
dhwtAROX+bYg7OxcQ1HxxkKTqA64xDxcYiehSGZBxfl29Ada40Z2di445DrJiwVnWD94KnfMZaGj
Vq9gVLwAJdyEB5rEM92pKmR7qYceremmhKoECJs227JUI++OvqpCtMuWpP8YH/Mmun3MoQVuJUos
mY0D41JAYQ9osxfMsnlhUWJSNFBDyao7+XSesvFdld3Ig3Utmo09ZK+Qt4PIPkIayHwwLKtJIW/Y
8In7TjBF3OZgDjk5M0xTMjBDcY12Oke8UBTFsa4c8D8oopkrdzt3KEIyIyVWj/7vXBdWqTHUCy1F
HE1S98T6IkBjN1QJ6tSfuiSaHG70lXZlZEQbX306f9aLgF/sIL4gnACllZDm1BAwOgFrMV5wO37q
kU5rcQb53Rqxx1Pq5Vy2DBe7bFnfluGm9NPdg/u2F6S6XmRagyqfzXR43+sXjr+V0nKq4K6aJMXG
vXHmOZARgEjpklcbREHe91WhdXFOex/hZRWpg8ufdMfTnNHNgN5GYMuc/2mtgNMHliOy3yhffUgJ
j3NUopSo/sDHCjO1i8Iu3jJN9LV+6+dUyhLpofpRjWOJpjLiKl3LEgoQ6NqhCY279Ty0LI+G8dE1
pWC8Fw7nEhcqNbsLqyLOvTW5AaLoZdc7DJgzm449SRIFBgkoHqdWanHUWEELxDgdWR6njn61KLFU
A4OuNQD3lzJo0jYILWmGlhHZf4jpeflvJvz/yAoIGxylazYMbnSTCNF2tmSQPICBIzbGDU1iO5JG
tLdgG66XRFvu/6AZo5nHAuhKav7Vc0n5zcsmkF4TTxMhJ6fP2mvL9vyPfXil0eDojbU2mejHdOm8
C4+gQaTwRay2IS7Wa2nOrARswoRgKwntyXxmALSUPliV1gPJgha0z8jv7AriPrwEdgDuxAXee3dx
xVbKz+gZro63dx03RBtKr0X+SBlHLxr9kvWNT9vqvbVcjb/WosilbG1EwbTPYxG8Kor2jtB6Vu2w
AyITDIjUD5BaMC1hEpKl4Sv3mqPvT0M1rhjdNay9DoVoFry4ygLxmu/eMXeu9sttbfxRYVN5kskZ
TScxnSkicGvaoFI75u9JofdgblZZ05sjqqIet94SyEAmnDxC3QpPNYNq6Pc/TryEg3Ik2vpFWxRb
S0X3+kpen4ARgEbB4q4QzWaD1xXYeTEed6gNCZvDWAd4jkBm48HwT5AkAoaLtN3N15iqwYn440G/
kj96tQUd2wAxV+NmkDNAFjlq0i117J6FudYY9khuMp13ibNCyFbzkkqy/WVCzwOuweREECyfAR+J
Y10Vd7ieWkrs4GCMxBkUc3lpbVJvQvc/63YSOC0eS8M8cKOxCZTV3quWvStrO+5fOTSVzznAMmqy
CEgqBOiIHj21yABPWbZZ1PQw9oHSYz0ke6yzw2KW81KVut2jKMcx1BIfaqn8YVrkNZGR9zWTV0Ed
5VO0E+fE3wevmUuRldBsy1qQNHSDIHRNH5W8P7mWSQQgBNdW4FGuo6aDvxy71kgX1+PfIDcsNNHP
3NIsWk6DoQBOE1vndn4FY2bjrKT22aVemu5Gn0khW/IBO3+90ATc+ICmh3q6t9ZnoD2/zYOMXgiO
CLdJ2iyDRMCIHfyWPdwL2KkOo79asGzuvnpXiAOPKpCbdiR2Xf3MR3atnpBzIC3izFY89+e6g/GS
cMfj6xkCKsFqMEfoljuMwKYFUBOuDLLl/9EV329mY2OafeFldBqVh1JXjxFXf8lMNrpU+IhXTYD/
j9g008wmmFs/cntVJJWe014/uFgUu8J4pESNUCfMNw3wMQRcK+d0K+vOHbfYUdVrIauD5phXPHnB
ps7QNI7rYVh3aV7ma0rRji3BoravdvoAxCykDv3GvooQupvCg5J8t24lEgXjp1IgLS8UyHWO1sS7
8ccTVsn/uFyLS9yI5uvzJOa/UQeVTEAoalH3reZq7cF1LoPsgDxXC3ev+toY0HRDe9h+6l9JXybS
UNNVcValIX5d8fRRK3im2Fa7KIxh8G1cjjgfjFl6Nqps5zvirIJgNagiJslsK6eVbsjC421iZB4z
73BhgpgjjYpIu9cKIzDbLo0LK8txXqCH+eOz/M1d7gj+nOH2EW6+Z2dAGWe2SMqagFXLSVtoQxxO
Z7DxXyjuRj669P8THzcbNHd4JjKmsU/tWJwEd9VPFX53dKwgcXsrOP6JGrlg6AOEMLbyMyfKNz5j
y0VVEBX+3q4h7hGnttzo7h+k2RufYvAIn4tWPJREhwDbAUnZo+pbTvfUPcaxwgkpMGuLp+e5FrNr
XwvI//sVQ+IQMSTXyUPoa+V7WZjTHAzHbUAamem3zbpr2pM/XyU1QkL4SGiTapPTkpHx8pxxp2B8
XJdSHO4/OMp4CX+CmBNXjN48k9dhygqPuA4xjgmmxr3UCfixqbdjtzCk2DEQk+c0YhaJBKmXtJpT
VL/nTW01/3Qf2e7IbPHKwZAVXVGzCUUSu6+CSe+dLbfoegcH59usImnjnKQiSJaszCJdbvxCx6qa
MYoBW9BgV5qcGRkfRZTlR5H8dQS01cRtByje/gbqG1K+qeDfS4djKUft8jpaHiI0pT/6Bsjy4cF2
6DJpJTexM4Q4s8kz9IeeRFbeeXmqsLLVve/ky+M0QQe7J2b7IKTjxfEZNSPgXc9jZ8ChmUmZyZCp
nFF/u78whNRpCuyQpsbOyfqMRa7jJTxWYmNemlluHKYF3ZCApit92jAHs8Q9wJy4mfDR/0+x8NMZ
0SvZTVpcSLLsgtqhc2t9oyEvYMMV1dYeywXyly2HoUH93rgA1LIPptRqcjnkopDeNZCxD7y0Ry8S
onzY8yHPaKZwPI8eGHZpacmJQAbhRGwWI+FZsjUQl7hpXcOE21g1nemDEtnK+4QS5+p3sm1CPMpp
+VB5VQ2qK6t+8kkavvOCRxLWGgQ04VnYWkj3wiTXS1rY4cGH7PMwU2g9csaIRY4bfECBAJvDMRqQ
XvqgtTuXfAiD2TyVBvBMlGSErQ4NWH9fjvZwW0NPykZC67RtFGq0qxYJtDJHJ3qq0r2yz1SafEjH
aGIQiHDnOmv8v0AlKI60p5i7GOhnwx5LiJQ35ufTTm8xOKei0wYxLUoVF8af2rUcNwUHtRE8GYK/
Bi35dx2FXSqBpVX/79f5fijyzTHXVidAG9bCvaGkSgMiRCqlx7BEf5rZn8pOGhizhoG7RAUzqA4g
2DP6MvAZVguy4GUKB+hnErg9cjSBoK5Crg5/rDEw7bzXYV2nXBwrYch7fuMvmcUETILRu0aF/eG5
efvfq3XJSN7xLiT/MlHEwr6jwFCFCbca01zXSU6Mk3vKlSBDmd4k1+L5CoThufWX8RQHOyVAbd1S
rs5rU1iLPnELynQJzyV62niQkmP/2JkQ0zuHHU+i/rTlCcak45GKuDY6CuqY08LD9mp859izgeMJ
e3nJ74FKHbV1CQey78iODCVLA9C+V4WuYkHHGGeIwC4EWSyfNI8aGCJPstFSXEp+7tmTYaH03xd8
zJaML0Vdh9KHO9Hqtm5dFyB3txe+FqY1EXj/1CVhB0AQ4TyQHF4EI5w658rNps2FPWUDwkvJVjv/
GOaZPM3067aMl/9y3rztVbOvspHELfVEFyUICmkxbJhTHa3eE4DQXhL5g2cgbbnoMev8zf2hYr2j
fp1/eUre6VsYxK/t+3IzykjwrBX2igt4u5Y24e/jr7Ev82RpbWcf+uALyz2myQzHjmIcOyF2xTeE
xeDTECc723HavrXRMCLqkrLA8mLEfa7K3Xdxv+aCp3zZyTqPn2D9iLRqLR0HONokszBpnF6PrUp9
8L01Kq36oYZ/6PREGJURdAYr0q/6vbP5x31m0K3TxqjukqPoNPcvLeBQ4gNmcEwATBqLbrZoNS3z
XR1uPwGG8dQfhnzUMN9oRih8YP6KRczQF6rwJbVuPk4EdZFSeMTmJUWGuHp173tZhfOZlXIJMkle
+dQBoI8BRKuO6hNADZqHlXs6Qrqm+3n63pDnRocqg/8+58yPNozQtgvrf1IKgTunusQS8uZyvblb
W3SOd+61gZ34a32yhK+E4HPYWsk5CeGrxYJNFFU8dOTsnoR5lP75lbAJzfoZh1JlU/WXVxeSLDeA
leebWx1gNrEl4nIxWzrnV3kup5ROLBVSZQqXgwBq+edKlUXVSQy5Q/MqitDquzKi46H3/7uV33Xn
r8v6+KzZufQNrFsPlZ3Di9cgjHLb4Ug080oK0UJoD3+Zeb2NvJs5E2KESomcJHCamv13i7A6a8to
34Kmo6BZ4FG8XsZkvHMK80O2mHXsJRLfWBBm1X2EzkKoVRRT+ZM1EuQBGMxeANIBiAsoyr5fQLwT
KQCT2deq5ZVdxX1eOhE7UT+9lAuQ3o0aLd8o5Ep6EcRR1sqBTgZoGgrv5KLHEry5xUwui1eG4lzQ
zoaNwS80W2Iy999SJhEdrVTm7Xw/X9LEmAL0UFvSGL4r+KyGeHG8RLWSTaXOIJC155wG6TLFNn6v
hs071HGsNq6qItKfwnOnD+ynP3ee9sp9lteONELYQkAghMx+Ep0fdlGJTRwso4UufEjZcBcl8ncE
Pc6db1Qaw01lSBgCI5FgP9tFqq1+DNsf3h39lGRHytr0Mtdc3fRmxHleH4niQWKKO+xlEnF+87n+
sufGEFr6xu7H0eCSksI8x9swDMt9r8g07d0Y/V7rzEMI/XF15NwkFk7goE+72CDKw+VBP7mdvZtL
BDnThgPJ47qk5jUwKTP/ZGPdSfmEMtO++06R0jGlbrcwJO+FhaPCeDkv+0pWD3lb1nyAbDFrvQ7r
jRa2AcPIaczu5DbQaCYcOTzvOzpwKn7w4DMuWImK0+c4zy+tublsS695i+J2ESAnxi5LTxKXLnNh
xFAqRZRPnz45I4YTmrdnHScvlUW472ry6p28rZjXwM2lcnU8XVlsOlv4GF1RD2qh1kB01iqyTlfr
Lv7f3X154QbUQ7jyg/X/9ZEH8XIbK0taLsQCrET1rgB+eCjjWKCEamqHHNrhHMgovRPnFVW6jsLU
wKRkJjcmLeB+/D0mLKRXKVp4JfLUt/mkGRJOP6Ku16iX/KQywxnmCQczq9LXd36khtflx18ChEf5
+4NxXn4z6eKQcrtARFInGTk2ex6n7fWkbMSApk8nH/7NPkgdlVc6c4Ed2pT/xT0AckCYaIaDKiWv
Ujj7wq63T352tVO2gG3OHtOTta69EzmleAYhdTXCpijd2j/cGHrYAca9I21E6ctcdeEJEAc0cv3Q
GUELidiqDrcXfo6ELI65JPR5D/QkXQf+fa81AAIOumPU+4L1Y3aDwUYPfaWAHQsQ2bp/sVs8Qt5P
AwVBjDXFb1K6Pdj01e62nu+02s1/MUV9btferFW+w1uG3D7/cu39KsLcZh1XQ0wkLbzdRoscJ9gK
FbFIO25uNK5k1oSf66eFRD/knHGx2XT1S2ZGPILlDaoyeLMu6V/ovdqYwOkbs6R/aCCLZSLCMFbo
SizDAEhwdttuS91RFhT65+jx6nbGlIYIwTO27FRwY8cLKNCQs9XfbapqkUTjXUctAVL+/EU4zRYU
zUirfpWNPyjSGwiQYTbKHQcR988isrIcQZySw/RZpymI2xoy2JQrjSUGmjRyRVSkF21sri+VzcAu
x+KEND8ls7rVdx4vE7XtnBgWPLkYxI2Sk9iCzxdzaTSRpfSI/MdjthW/7bHbYeo0NDPihcZynKGL
uavCSeXg/ihNeATYP8GCk8cKWN9PD5082Gvk9cqulKkD5qNESmiVTiCssL/uignsK9xzfnJOJcj2
IJHxdQKzITGRZymg9bcTdiNBb8SsaIQGJ+XCrVxpDN7X8RmocFxB/qd7UlTbWYFr1iqX5qDpMoNB
2k64XZlFkMk6X0vGspn1/uUa5TNrGtxEQWM2S390nHRWIuh3JpMdOpAjVNULcPtGzTbQwsTpd+ui
M0JpwwLp7J0lNw1YUK7Am8hwiW02Zlpvv8OAsIJZHsZ91AmWP0xCoLvNtzlJGZhngo9tNhb9I8ty
zpJZRl1o4VIew1dmPMr0vc2ZYP8mq2BS6DiFmUG81C/nu4FRuXpJ2f2bZoT+WPkxCa/YPlRz8CgU
uXytzxxtq2kM2uh0DMqtJMbcWOqtv2uZDtYj9OPPLnLyo6xe2vhHwnmm8ezMEL87ZtWvGSvXLrP3
gK7tj4FKPNeQ4t044A5tjRyapSz+CWh7hKKCJFrJJ/zI/U8YHvUhRt99yvSlJJj+4sM5JYqh7U64
B3hyRmHC3GZNI0yCjKWKXwbaGjaDoDT9AXn14+mvgIpqzvckYISbr0XTtzdotuDZjoVCDQ/WQTsj
NLdc6ws+061g3vZajqTDGOY55vL4ba2KnWsa0Q3Ae0uI59c2IyAC+8T0TUYKJ8gA7OUUIEE153fm
IB8CX655a/9HwpaHOnDYM/Fs1onlVr5zjkxsV/k0rKWZjV6msk8n4upW89rvHRxMTUgIXbXqLg0R
APQPDgrQfO7rwZJA4BhW3FkO9QUZIn6oULswWmYlX7ZWSGROXHIXYlMjRSKLZb0H4QldklQeCuTM
nRbNI1ysInQdtJG+dzzkVAeLWNJ3JCjOr0HqLbam+84s59M9w5x62vIfMdPedHoHbSn4Qkyn6wSO
j4x0BTToNyH/I3boMt9W2eVB6tZ9oapAg/6XC+78i4yyNgXEoXelsYGSidjwAbZyZ7kKLo0gMMvN
MsU3Aa2PkC7TfBGMOY+ro20EbMrdkEHZiYxJFurfSEGBo1gjb33Ky2ak7eNdHEuSDwVZTbGb8IXf
B91OAbclrxQrS6L03/iH1uYni6P+ec0/FbOG58Gz0hYcOh+WpYDMjvQyI3vYVVlME1DpmsvwBpUq
puJIK3gCi13w8/cjRXw+AqR4GGOeOAgRiwa2GU4gDVWYDB+XB74qvGuXN2dX+Cf2GmPnYJQkqU/3
MUCJ1ktDxDwrEaS2UlQ5FI4E7lh6QM7B9EWTyXNm5aH2XKHyHxBbtgcNzra6JGiDSqsfbJeDtSgp
mAD3Wnf5nvTGz7CJZ4vJhSguMK9WRCFvmjuH8VewPPa3FMeGJR6KwBz274CoWJ/R8iYV4ZZf0SZr
kdMn7GjQ9ZLF9xYuXpzxfT8FmHzwZTZSRi7tSHmPz3V+QE18p85kJAmr8Ycku9OzVz8KZDMy3REZ
2gpUw9F9jqmbucnjHTjxhKmytyLAHpKspfroZjMnro0p36w1RNBXCR3zU3duj+aajmqVkHWkWIfz
Sqz57+5w7WU/XDB6rXiaVg9coLgqyvKUNoSiiKgjy9RUxxpEOV1iixSI+1UftPy4n8NXwwzZidKL
srBNJHirs04lzMfDyTxXVOcKS8HHA2L0YnD3dwKysBBorDKCO+vhB2sBAfpmoe2nzoOaL2ChIy9Q
1RSryNrdHMF1jpaENPsgMTv548gfw9a+SdeqHnA8u6y6gNAgrBljrm7f54ETxLaXfjfJ5x0MXNZm
YRSf9D82rebe8StSc9+mGRKowRtGusZLRW7Ii+HJN661UScSB6GVk2n5JgfIdSpsbM3v4Hpiem6r
sfw5dJxecpY3luW0pmr2foq6ceS0ZGOaz2htkbvQBGLL8OatRkS0tzKzKJ5lT3i4KNEQ2IgUfwWL
i69w2vmM2FX2TNqYgSUZlMEgQ7UEDY2UVLZFK5n50hexEL5XG2/VMVa36/w35JRKe8R5rmP3XFFs
1qHys/pP2FAKL0z2n2ZRSKJWOYcIaZ/9bbZfWVN6VKWTbFqJM14n8IUyzEWbaHDFzRgxl0SA+eek
u3d8UY5JiAz7b7LY0YvTx6e4V/m4SgYLq+LibopcGoWmHcYGrA4wHhAGIK46XyFbTo1mgC+aPxm0
wOq4RDvqgizeBaufr9jgxTP74zf6lpgOOjnfdDViRNMuTRzYg59Q2GiNclATkrf3XMShmpO+N8kX
arKTk0WM3A7s0H3BzL6JLKgtnnBQSRDVHlLhjunaivYWIu9YhPQVqqecWgmQCnqjXV4Y84Nmq4HY
g9LLPUbf5eV6L1TLaZW0DrHIlgLwCqIZTIetzh8Mz9MKcgX+9J9GLiaCsXX0B3bwR/AelAd9g2QR
HgeljRhzndYG3uQ96nxvtLNmUk6/w4JxonkjL8ugEuabXlWkcyNcZ/7ZbzxLpzw7nmZQfFiWq5vE
pxlBTgGnY6vjNufl227eWFHcQXu1gfuEClx390fqgakKyJGpWsOZwcu1LbGl5K/AewdnMO4hq2IG
qepOwfKuIVpvMwVs/1dANfwsP7JVUoAHoVyCJVkUZabLR3bSmVFQNd2l8w+QTr7AdFy8E5ss1e6l
K3VdMu+uuLgFcZEgr6p4Pe4WS9/Bz2GatZFuUIzbEGOvyB/s5RsZBkhh+9psraJYk4NLSnXs90BR
nbY4+LsLHn2FUsE/VV+vMW+/sDiQXgiearsS2O9I+MJdBHMKHnOpgBluVUx1+xyVwZRFW0S0eWGx
P61EXi5Fck8hdeH2nRxSetOoHHPfW8etHMJIGKOzliOZqGoGzkP+aStldSgRQSMCF6rbWGof8VX5
rzzDKxSZ1NaHTRBMsqWGm58vUtWkBRkyf0qanBT2EU+KCPUKSlEM2sU15hkUaMlsh6nvyh16saXl
42R9y+IHzYPiOCOy86qn/P5iDxImCILqHG777oBVIdQWjb5c61bkMGDy+7ZKDozGI2D+QbgUuRb5
RPke57s9XoC781/3Yg/4t5P0G0EW4DKLfUN2F2pzOiW7J+Y/RMwSHO5xiA7uFrgQbDf6xvY3tLaj
mBFO+p3F4ctKDkPf363zrRovCAZr8USdBH34oML7vrNUdN+AD5TfbZJEjhLdp5HRqWdOUSju0mb6
ix3ohom09b4EMrcig/66EQCPiWyF9VpNIE5zVFOsyLJaNynzwqsEAo6LoPxmsLM2s65QOF+/k1ii
nGfJEiu2+utlnJ4qMW1l89oL7BVQCCfznVoqafD38U5XIRWSvQutofMZ5qLAIlsdW56CPa9Nyaud
p1Fwn6UtFSGBGx5AkY6yaGKgMU0qox9Iay7O37c/vt7xZTW0PbXzP/EMiPAcMGIU6JtFJrqfTPTa
GewIp+93/KfTLVvMVp6UYI46g8C4MrYgH8OnNI9OVfr0F6Bqy61qKx4pHhqdqscyH/8Sc6jr+FGg
IiFdyIKdMlzGsbhNQebA8yODOiehDOf/DvVoEwMhSzh6H/8mzZuoiU6KixXtDy0+x3akLBE/Y28z
hSxKiYSfwCJ5R1cH6nd0NKA3IkTTP/pKmsAnpeXipctGIPNRGN+pZQ5Gx8j6xlKXYXW2ShHztMH9
cBEACf3UgiIkd4fkfuCwKxqS/wJhzYMKrY5jkL1mr2nzPmVMtG3ETsszDU5ICk+/UIH8MpgKfb3v
rjn2Gz+Ca/01FbENhsEVi47ZVWJJ0pQTn5HUIRwkbyTB5462rWMuj8BmaRr7SDFR5Y4NN8BUzJUK
91bLlG85p9WGG+chhXaX/x4FcJlQxvAiwZuxUoz/hbgv59L/HUdvFx1qcmOFTixFujEnnk+byQ6E
YPYF7OVF86wt2IVDBQS21r/woQZPrnQdiGCA05gfn4vLuMQqaYfN76uTQL9PRuCIENVf98eSop4x
c5bPuAMAPMHTlBnv36YWrRAs+N3xwVS1TUIdN+5uj6mawiOcZHWAIbaW5cWEb81k168zxcumc2ns
EdzlPADF3PPBVvgj7TdullUWXqVkahWoX+2+iVGdXQWlUqa8awn1GoUXUCq1Ep9/9amqKbwkcMPd
liBGfUTzW1c7J94ep04f+Ry5rW31sWJF0IlG2Ekd8odCCgMdX2Slvld5HPvX63hiQnzcFSqB25EM
L57rOp1RkBS184Xala50LLZv0ffmgC9Mhyc/Z6XXVTPoAON/NJc+0pm4SEuWRdKSTHHdwoFO1gUA
KOGzy1KVCJ5m+o7gY0Y9AzQQ559gii6NNsCxWa8cR2lxToMJtluJZWeFSWB5xUDEZxz6PFEMnJXy
425UEByvCcYxmC7z5Opl9xwJ79effXw2lKiA5qSTxKhvQfzIFqKPsXsBvLxWsyuT2PRY5ZDG85Pq
5uuDwE6Y1+X4QnI1/Dg57tbgjpil2pQzyWxd9VVp3o9h27NEod/aTKdz/kLQVWtvW3Zoz8RFaCJM
xRHrL+uyVkJsed5KefJC+cZKPgeiyAfqkoJRuRrkviBGvntTXmRx+uw4HBeO6PD7SUh99s38G9pX
6MsPKwIeOWE5EUSxWYEDHTm4HhLszsarRKshCDuwCwmqA0ly27YNDNiUbdu5MyBu2wFRCp+e4ZFX
0VjsjIgOT/wUKhPmCj3TttbgFO2v1O1aWuYyQY612Bdq5dprInZf0bDMRFoP5HexyBsOIWxjWPR+
o5VZb1LUuEHLptgEqbdPiFTgHS6ShETbqNnHk/TN9EpBKDGvadAU3Cqxp4ZWTXCkrd1m/cQ2Ym68
3a1+nVzko0/rSCluRHjt3mjhsRe9nHaRDdDHeZmlZ9RSP2AnkukysfbMt+h/i1nTRgdlcaieAjWa
f4IRTGxscXTjqyb63DBisMBL69hAkYZgCqoWQID0yFcIMZzPH8YGbk8S9HfhE+5w61Cz2ekEoRwh
eKH9tCslbUaBgam1/OQ2yWomAjSIowjyQef4mKt9m/Ql46WQ2goMec5IViHfyh5dgrgpC17sjUFk
BfnhtA0UFqxScilEmdumj8jGPt5sZtX+FCzhNPypC/dlgl0PEQyrV7BfOli8d7Q+Jau7EidodxiW
93FtxR6zj1UNCnOzEGPzFKy/1hU7defjXzEDmvNlTVUrTZ7HzTcE+B0tQbUaR9ZlLoJ78e6xvUjy
vONIeS1bc1sWR+6wINI51krsD6NQJ62n3ElOzqs0AZ2lMeOG0cxv/jTyVu1iAwyW8tGN5+FRWnFH
NXbXV5Sl2IDWJHkN0aQgZVgqBT8kn3rZkAHCjB5Lw8m4KyjSxaFAN+Qs6h6UHaABbvdSb9Zurq8j
Rgz08qAo3gp8PEQAL8hMBSDGHeyPqcqVdUoTkn5S6tlkXGfm6zuKMnd8joPwIxG9p84peSuj4qg/
JVptvFP9C6YzTtLs54GDLEleQGTdFSIRJeCyS36r4WUjrQdIUf7dyUuGPnZOk7TB6DtSj92VuKii
EOaoPaCjZiWFFJycb5QZkdZFvKqO3TIzVwOiNo9KLqHy/kpAy6ZnXxTxWs+mfrCAv/JxkYUUd8x8
vh8WOV4lVJtxb5byZ0jbHNLrxRW5z4QzPbHwEmmENDVwQuVkeNLWywsdCkDbAX2Em6mYYBExaTBw
S7jgrgqBh27N8RgW3+xInYDTCdBaShxKU5xSWzDCw/knfzTVuWFB+IFUmv/PpyQljOKDTmnLSQt1
ioXPobwd8E77LhQKE1LFQOQeCgHOeWj0aTcU37z1aHUBCUe4vj9oAdsmp6JXwMw9BY/znG6RQhC5
ATH8RSKmzjKkAs1TDNM8x+uNOevmLzo0s0kHaWB/Ryv3jrqVJ7dyulD5L3zCTHRRuLtxyGcTZrkZ
ypoOBROz19xdEmLjtR6RStSJtZIRleDSSLga7QkeJumRm3T36hOtExwQaer8PuamAJq0wym3vbuY
YiPqSI0F5zFxjM5lHcXPSpsQrJ7o9hXa9SuolFVGpOGZIxcZFDY0LJghKwUzVpf0h1mN9YhdNbJZ
ZVM/KDqrqYm+UfaSbN26zYKdnkwjla21nalK71OTFDTuAA0toRqmJD3XWxdJ1dh/3AyPTUKHRdXB
apFEZrBZHT00E2kC2uQCja5OKuTRX7dpzxQRFFbUqfXw261GPv1gtDkIRsY+oKq1OGy264Nick0W
e3t0uSX4VLk0jEiNkSUMqH+qZ40BmGpjEGFjXkZq8bu75oPRq+v5vhENBhdPOenWwtV/AFdl+oEm
5lAgTI8v2L08/zpf/i1wTi8m4qSXEgWtrFcqyDPyoxqSP0zCVgYg7YTz//ts2umYpHxNrpkPfyzG
tLHZnTZ40TVowb3JtdCLF8pbqMx2nVdTZr6WPgH0C3Z+7dt+KbCheni0kBsB1Peljs1tSlEXXmO/
VomuRrBIrZhgXPZZgGwWJrUqpy9BJMId+cWp0/1G0RrSZqeHVZkFmfhN7xuOKHx1vdTOkNSYHmC6
tN2vgGaozuzWN7/y9y5izgqs5CYu1SWGHwW0EEssbGeL+3OEMLo1srKPhpl/NkYM5gXS03ziQm+/
9GbpY0eeo8n/PRqhBBz3orkQu1Dmge1llKMiuIab2DZhEWszbppachRUQLnFgfc0TfvbhzCJM0UT
Ieyd5LJyxYoV5pXLqBvWyif/6xZr8rtSBRC+6+VM0jv4m7bOuHT1qObKB72kb7KYN8HhkwJSsech
ahxV6dsn94yc7TIvUzZ4qDS8L8ZE37Pd5zR74bwfD3YYZ/adm71bn/3sPQafAqtX/JTFMcXDxFBV
jnx339HqCL4b7lblm8EOJqJWTN86ifszBJQpHA1wVn5O5xmhQHREagG0+u5gRTJZ/nZugtLerK1v
eBjmYqtjmJDLuCDs4qZUdKkLnqoSL1q+tajAZMlZWIxP0BdhnlVvPfSqSOrHTAE1sNovJnbyHCPB
xzBSDOFndGCCuACNIiCgfFbeqJmB4HJD0wtIWOqw8GFopu5tASSpu9RZo6CfsXOf+KRst57ZQ6QT
5jfbUx7643pS267Qq5jq1ly/JVU7naDhlBrQ2GiEEnrlja77G3eAZWb2ABtJFxvCExRGSG/clY+t
xyL6bJQPOERnmPqhVgwR1MGCRmslcmD1bMPGTOHp7+y4InJ3uCak/XDEqmKeAw9YPRlbamVUoYXI
sbgzpq4HeadpkHjamChnW1E4mJIga4RKcLWdOxp2j1EfQcp537v80GBCkG2o0VPYHMVBBROl0qGR
5+mrDQi2w68KruF2yQzv4iwSdqxRZ8Q4ZRFYCL5vJP11o4OMK4axhjy/VcflRB9OohURBhTafaNS
beuSuoPRd8KQL9+JAIFSttIGo8YUzIpqnZoDP8Pt6juMLNrRsa5t0Sv/ulghLsm5m+aTDOYz/DyI
nVuP1CPXsjLSqE2pw8alcBzo0i1GPX4NDU8g4mNemr0fgagxja26hCQLGeuAPcE1lcGpdQLvVAcU
nxublugLaKbMiiEDd0gYXfOfgXr67wyBd2pnnuNDi2SIfbSZ6aaaEZmlHFe7P8s8ow+zVNuGh+5q
MYnj7som4IB6DF1Y+tYFEE5oCKuNb7BpuUpE5tTGzEAjZW7n4R2ajjh3XPSl0DaccMbPpp4pd3E1
C2Dqs73jFEZnF4CevUTNxBUigXKErMCBVoYOqoIoJ8UVQlaDk9W9ZHqCAv74Q3AoofUwh5B5qrnF
Dfj0DfJODOz3VUjvu/cGxOwDcVEQ8gGP290+9B5KzzNvlM2DccX0wGwUU8vL+e4VeMmQPLUZUcxj
7/Yhu56vg9KApv269IBFgIbEZUm0l2/RJ9t5sf4HxY5BvzIhBPOH4cgivjqMbvyDNpG2ZH9ie5Dz
izoMB9Ic47vLkGeajwWLt+PsSJd2wC+gAfh8Mx20xF3oiA6ykuGR5bY5ivDMLfSjYR+WDDTNo6hO
+NmVoANmA4pDCf6txdeYWExm7rL0tE905yUxyXFKq+rqONLvezb9of6upWF9JYkydF3519RQJSKd
UsqpzwKOjHKbUPiAlanctJe0Lg3A8eNNEeiJgVK9n/4tjyKUC3hb1B1ljGaIg6rbd1m/CDMUV6hS
aNmgQP7uL2vnzbYUCFV94WNXepl+85yFpWTZE+VqyUM9OUI6WNNevC6Dlli7cwvoOYHyO6gFqrkk
48sSRJrWPJPbArpK/T4O7+sNZndEHUqsYpVWsIqtAPXU26PdSS3OqafgRM5OhQWRhR0bLzpYBZAU
ideVoqwJXBt8k11ZCyQFtEGZLDUv9UGZDUaypEr/SnKvMKWpTuNUwlXIDKvIG4eBwxZcyLUvilmF
F0EQW1JKjLgUCItm3W5tVQZ1+QStU4+vCIlxmIPxq+mNvR3WZ5vFPnxFToR5azZZ3ab63Z5RbtV1
uIJsxWSrrDMxvYa2FF8+i387L9jYtarTPvio7lwM3shN+T3VhdrhHy73vh8t+bUvGdHcJQ47mMAy
HTKszq8wjzUcli2vbro752no2kp/WTJFtS5kHPQyJjKThOk2hNX3V3LaGDF9pvT+huQLlndoybI7
RfECAq9WGoR2fV2Fq0WuiFnMidbEu/pDOZHT/aVHQAk3ubgGCP4RHZLQDHcaRVze2dHHXbBb9R4E
xzrPL2UkeEnBa4Je+APj/H0eqbJzfbnKYRURaAiy53VUPn79/RnyKJ9QDC7DBEhiYIhBoMkZgjy0
Qu8E/D3eyso19ogyPxusQK+WTjOFeeHDKykww4OCrhjBejf+7jtccO/SzuGd8T2/017Zs3trJH1C
PVhvTIZcniSh6BkbzEUpJk9Z9Qu7rlzUWpQN4m5qAXns7hkefoDyvt58SyIRoRdc2elcTu7ptBbX
m7bsfxS4rRJQuqC/DldpuT0CkNd/GkFtJnJuailGtN6hAEwGLYgNu4cR386SGxoOb3JM5A7mcT+K
u9BU6+1Fj/CCCZ3xc9w26N9VBoNmC0H3UjLeNLF5LJLIUk9CFg/mEjZk7b80JgCfbnNV8B52qrOx
gwsyZnWQ+5EWsSJR3WSHx4pFbOTSl1RlP7rfqaH64MX30izShe6Ue9KUzunq8FZqekeA2dr5f12H
SCJPC0TcdFyPPtsX5e9I+v/GG5Krov+xM2DWDSnN3y4HqWRpWDYiEKGscOO4CZVjJ8mcUxq2yGXn
sR0q+ZM/TzJWNb9GPHBK9sByD1SKPeKVZHDdpFZNl1Xg/7/IBDVfGgwh6YLZAyy35g+eqc2B0Opw
mnJs0eKvdgxVN+vfe0QW9nM8gfQ7LEhbJGmGIWpY5jhdUX9Fm+kIT5X6pjrmjS5sfhl9Tu7CBUC6
kntYtM1iwY9v5xB0ZLXfyyQsZTm9OVp3UrNXMKv+6j4dl0mQKA9Smcd1Y2zuAxHT8fN+S0+AwJBj
HCJZYBKwEiurT2ViWqLGyUxOCiDDZ8u7RNrhuO+PJRyvsxcmFjC/Z81Q7/Rbb8afLWhpbtkYYylV
9rLIXuQp57Fm7ANoTXvygYibt9ljTfkFiRg0pFNfqMOVKIn+6dCj/nBmofj2eRU7S0qf+Fcs/2NY
ZlOR6HUv/oHKE9NgNTva1J2enaruyg32jMQgZyoPhgjphjZ+Bf+o0U2dr67QIQ5v4Onjhu4Za/XG
hh4g5riF4Hombc0sg/yRfbACnttzCdnyqz/4IgiHbZjGg0axPNjZDQGasKIFyOEwec8uD2it0FzQ
MJu8AepzQmYBAxYdm75NmfgdjtHMQV8n3MxIUFyYJkv3Jy5yV9yJYK6D1Fswv2GOvqpVAwwv4Wfw
oZkkZLN/7OJk4lGQclnGEf58MFW417Fc3kZCV1z/T/OyjRUIgSfUtiheVZ0yoNrcjXxV8QeQrzf9
fscKNsD88y2BS9MESbBVFr/oNyCtWqeDwP+m7OwKcqEzeuO7I97Jt9Buy2EuF9pZEdPSk4qf5yVV
+z8U2mCJDih8OT5A2C0uFv3oUKFWTvUBPezPOvDqyvccqFbmTT0hAkjQwHEnpHCOgk5hSxVzG6Rk
gKNBFH4E0h60cv70v2iRFd/e6Q+bGAsN+H8RM2qCV/wBd3lJ3oYnOg4rwPnMbsyoXDgFLy7y5p06
FK8wPt3gZ2tp+0aZs7wYGekLvgL0k3hBdsV75+pHp+pk6Upxm1QQlXiwLqirRI/8gIz0f+zC306b
YmOW+9rvqWvV4cNWcM3Om0qFO8NOZLTpOezkky6y6Jj1GyS9JaMHc4tosSiI84cyWD/MNbqn/Q19
l/L5QEhdIj8CcGoxa4CxN9TVQpXFQhkPzGEJQw6RNnX78bBEyLThCuXh3Mr3k9xMihUIeC874t+o
GEzggDDhX9h0SdKU5lmvOiIJPPTlaW0KuFyUiKHrUUTEyGJemDZ0jYAGGodeQJcZ4pUxryb5fM59
iRBkh2a4c8tD65mI4gB4RFRgXqDx2u0uPMeHa4OwqJqjhHKSOA3zBN+n2Xk70UjuDik+6BntT+Xo
kKuHvDL5GH8eOgdLmDsvqCWuWcOgca/kLwTkZJW+QzUk5jqW07vlkNtE+PVRfjJNA/zvVjsY9qWa
B1udugfFR4bquwnENsM6JoqJdREzFGDw2yZXLNhzRadOAuCYABIDTVOF8UGpuO0kqG5CC8bcO5R2
uYdCo5S+i/PsxtcSrZYCxpMiFf1tIohwNVdDnWjU8TPHL1xcjTSuCYWKc/W37oW8bOLHyTBZhHGd
PmHHelxk6Jc+bCR70BZ24beWjO8zc2daFMHjOdoPyUrIefw49wJEaVf/Fs7fNY0xJ03QJfYwO7ha
FuWovbWhLbXKLnyzauAJUCcvtZgZC/Mhe9I9WCCIiUiDAmkryeH580rBsctYWK8+yK+qNcikGDOQ
gUlaBFd2iQUEOfeC/SpGBs8MFl0uwjfE5xV9wBBw5L+XHFwUzODJcwc6EhUC1lGo7t9MF6EAZlIK
R+qY1nxBRUh6xtwUcp5h6zxjoKXygXvoebBG+A7Vh5IX+y+GCsTDe+6AO7/pgy6+yIHuoqAIN+gT
3WTiTduHsave1Y5DreAB7U/Htwhmll0hZPKvFw1lO7dioGPSi8JIehPWKofNcPpYscWdliDOOX14
j73eug2gBHM6KlFmObgwfma3YXmTrQD1Vd9chH2kZbBvvESUmlcSWFdH+UxkkBPLa0qco0Oxp1M6
zRjgbligRlqGXfzYB4diQQDjmrXx/J/5fT8S/VfkP4Ey/Sao7uNzxssfCR09jbZZlmuWICz5HMhD
1ac5vbENZ4TNxkUlwoSe1P5ShXhmo23M29y9xTvUMN3hSr96qdpfZJ7kRrF+102azeTB9MsliPzj
UliV7ux9quURbRTsSwj11MWhChkUJzqDpt9s2fGStUKPI5W71CX1E3wgrkZ0tuz06vGSJk39DfqV
O4EyKPO3X/B1Ol/dBBPxU8CzlnixARQYLRgq02ygRrVmagC34Zv61cwThm+ToIjmjAgQ9lryFx7Y
z3iGSOq7FgzjzlZP+Jbv+uGSGjHgdzFFxdpS/2odjodMKw1VhmCUARBrAN/3IBuLsCaZXQgTYOvD
DyEuvy6qyUigRig8I1Jr2t6BZUWAUEFa04UBcq6g9hmBeeUbKxf2eNVU4jiTYNsq0cadx+Rr11sB
1gEqdw/LpykF6LLGujd2umRNI/MUlwTY4+GEX1kqPuvAuMNM72TRAnu98uJMcPtD5OyseAc1PBPe
ojV9bI/vXfTi7ieiQcOkoPdC6nDwo/PeArDpyG5XBEMUN5kHP45jMEgX8c0r5oDHqUmhAFG+E8tW
iopbIrEUI/bFSovDnQIgiCAvs9ZA97EuSSbe0s55k3ubJ247iYrU8HcynhDOvvEJn/Egz9dwbWId
l5gW2e8tiob4PH9cX1ltgKVHEsAtY2tjpEChb4hsPj7orRwsQc3IsxIUC3yc40ohIWz5PrCKakzX
+p7CqsacbjgOlugtzjUD3AUMh4lVK+MdOPQjVd1ksu/P9eKLMXtMTel8Dudfwak1ioahJ+xEMRJn
lhbagZPrRy1RA+GRn2hvdMUEHXJYy41DIy4dbS3Cvs6g5DkcIQlCz8vE5zvUYLL66dydLrXippgO
Sc63+8aH8rNdOOKbZ+1eMo9U9MJUU/P6HEbp+/lHqwIXUya3F7SZuWJvkbge4a+TleSMvCp6RDfg
HwH69brD3lvd8J/k2Nx1cjeM89haZWFfesytxMALsTm0AINql4PXMFD0XfFblC1+y4KJYb6CIJ/t
qodO/2sES4KK/FhUz3TyX0Jpl3Jd4ZA2Uz0VPc37winfFnhPUiPbJc+D22CrcXsinbQhmPSyUrua
SdQMrF1E3QKYsgMPQfIKQJFlr0zHlJC1IyTUD75CUxbWVTyKXu8NhgsQkpHLsWJajZ5QVSjJ8/Z8
rQM9eN8cVHxQxaInsmaQ4g8aoS18D+FqNUNX9H7AOvY1smsyW05M4tS4HE0c2x1g2kyQAtpHMaCp
xIq+OvNnxNyLyZHF3uhl0w53nQPzHiWdpotKC2TtA3A8OXWFYWifSpVAZvnmxKFQEXfhdG67t+WM
eHDQm+Vdu8ucJGpt7tL2LQqVepUSrLQbG2l1Lf5gtTi060bfv/asOqFo3Jib9Fa+4fE+LKB6+I9m
kdHeDxSZ54b/G2UGQVJyGV8z7jB7uQdTZMl1kJ0zWc0RL9fwM+wrAjTXNvwNRIUGLg5ZCm9z0TZ1
clL+4P8kQMKor+jXbD5ncwwYhwL8hk1d8+IYENNiSGDuzVSnZG+VdSkeDj881OnCOb1IeG1o8psw
X8o5bk6RstFwrdOGhaFEoOHwPjrPt0LHD8Ljvf8/3js1gv5SJ4B55I+EKOrS2r8LUbuS5IChUzF5
eBYPoVdxhlDuQN3YARloQzrW0u50LuahZLCxTuDNmG1XnbXL1YXRbDFAv8zD2AcClkGlL3QIA3pw
HB41nn9HR8xz0YAnruLcUfpcZCbIDwo4ORa+ofLGeNqwuPpl4ILag0wZTtFyttOeuYLWTo9s0VhO
12/RGON8JxNIhABJwGb9G5DrQzSgSauqeyNRszcei1lv1FOG4wdQurdCHFsxn6f8VtW4QIivOFzS
jJRESk4FMUDRN4DVU2aj/CRa4ef+DEVTyJfGuDomAmYkg12gyVMSeCuT1Ab9NCKEHGgNJPf3IcjQ
lbbpS9mWMwsyITRz8QqcIrKD5U6rC753/1HLuZveFH9pXZmkQFGUuX/akpiIdyf8XxF9E7SkivaH
fZ0cLlyvzPc5IbbGsxoyCQEHF18DCVeyQEDKUvfwiiiyU5oMUz4gPM+l+ov8nvIZ6Noy2/M65FCE
VdLa4LpSBfUDUES2bImqW2tieZgNwnnGeLf1Yr3KaciVSeikyguUeA1OhX9BUVXGsLrb6VaXWpHZ
oH000k9MApnsqmll+ZkxhXTCX3/EPaRSmeMmAB33ZUpW2ZwllUlhP+0lFjobKYln9d4NIbGpL4mm
z/PAR8rfYugwdIjl6Nm78h8Xo1lsOBLZzRTdBrLPUP5gXVVS1kBDFJfTT3OhL8l66u48V3++QchR
Lq1v7TL2WBWsErzLiisjk7NZbB1UqDL4aFJQLBLdblmSZoGk35i20tOsTY7ZRnnEmYYxJ6WGHA+c
fH4FQnFtoS1U/W6WJvoFTfXWhpI62vf083MW4ZIBJXpPMH4Li7s9JMrDewTx2HdB/tJ5xd6odOit
6JpvItvKv24oiUfPc6UoTUEsuRbqI1jLSTqFbAUK3WTmIMH9J8QwxJTanzfe/SFr+TYk7oSoqnlv
ys3m4LoW08kR+3v+eVgRBW2SwdLmdUiMPBmhnGnNo3+e2M1G8/1KleXtNfeXW+EJi5Sff7/iTSJ8
8rRTf6fqpnZUj61UjdoEucfMv+eyJPfOOcLT1ETDM53mT+IwJK8lRO3mv0caq2bfeEMsZke6bCEY
DTeTDC1hQ9UOywpoUcqW2CDft+T9BnGKRZ2BWZ4QISwXWfrELq94hf+f32WghylIBQhblSSrhDIw
MHGtmIRQxHoTCPko9VjGnDb3RTFn6cDrG3fMroTHbYTRbErFImirVypK2/mpns++e0Gzp0gyJIQg
DxXjbW9cZkKX2hv47glcgLuPpduLjcFbgRHDjHfOVBT0qNs269iWbBHZOotVgmk5gqiUkXWkqO1k
KgSSq5lrSf8JUWNnpK2ZS4R1G35RvN0xct8Zx2J2dHjLABYr4yaPJg8ybRQMaOZfAVDVVHGjOjMF
TP8H/EyOlmtzzyV/3u6YUi55s/yonLnluWFpIxox+LvbbOVcu7qcteEhhKWzv5lQhimGPeuG9Fk8
QN4mCgJ9wIheN1j2CaZEed5GAeCRRye5FWPl2Wh2ijdQTbKcSbQNzaI8zoYgok683aciakO6f2zK
7I5EmwexR96boATWrYGqrqRM0nn73Tz0aJz0J/hq2+cOq8b4MJeBBtOMGuwauzsNxlubIyC/QkTe
yQaRQNhN74W3BXQPzS/+bIF+8p/bbnyua+b+jF2obXcgXTbd/J4d/wa8+rrDkh3S1OVAUXRm/8aC
I4e0K0dA2lMgZrE3AzdlDe5ONB6gfa4hh/hRzR03WO7OK95bnZVkKcHlIR3mb4NNXOIc2g1G8B6P
N/BTwQHTYED89KYX1BWALP1oQ/leqaCFHDz3QpHtvUebOS7inCsrx68jv158ewGODRu+1r7PwpH8
Uep4D8CpdLepkC8e+7fmKuZxX9J9STtxs5tiVHnPd4px0GoGEAFDB2tdgHrDNA2p+6qkNQnVm4Tf
UfXekQU+i6WU+l0rPU15IolTf2va45mOB0VEu+jZl2EEZzfT1tyWonJHJFIhz5rvmt/kOydiTErs
A/YKiJ1kXDLkA+kitWriVPYbd68xZ4vfZ3EVqCYbbrNNhMj4f/agLqpTOAWeqOXjUO7ojJK00p3e
tNLMrjZnWAUgSO+gTc1MZ4AfzHsyLvxD6AGL8e4C/MZ4mdy9i3DMHSJio8dRXcSzSDaJe4fO4uZc
BqvWmFTxJ0XBAe09X5BOWOeXWnrWA9SOjdLC8rmo+JsN2u+v6Me5AC1w8W3xbk7ormgvtKjBopOQ
2wydznv/v6R/Fno4/87+eV3djEoFYtUQKQ6nYWBHUy2q34KpasX1bs4i6xkMjB8qFzQDcmzyEAZz
W2dRD+iQOR52sWRHopo/Mi49b/AkT7Tq3WjwHOa/ebjoNRiN5NYFUsBbVxvMHniYrYUP2G7qGimU
F+CJoABi0CkK7QVJk+8Zgb/qhhi8yU/DC9F8c6hNwuym49bCMMtc1IdqCfN81DXRVILDFev0vls4
K9K0W4QVvJkrgx0qNNMWcbZqBRSBRS8hxYnqcT/Q1q7pyNtWfDv2CToZ+JWyJCq58CHu3TOd4TqJ
khokF7FzEBmjfqYz4uyYQiCq50R6W5TGesqeIx8y3/p+b9InZKtDCD+U7dmbdNg9WzQIhGUs9yb0
8YkyCSrvrkBEQW9K/qrZFvrsEpKsrLKVmkZu7kOFUhK3xzAseDn6nGoK3o3vDx1608X4SvYqp1aO
qEhvdCg+jFOD7hXQGHRD5Vu1D3BlfurXIFjgJXLJA7ZatEp8EdtLqJRpbVjT06Es3UQPPMD+viuI
f1Qaemdac8JrjgWHsdb36lk7JP+So/OYir9lGrnrXGyzFzctuNNBYDKFHRUhH441Ok8bKHlaMyKE
MTciEm+nk9JQJ3WwWRkvK7ewaxu/GU2uOFnI7WFdC/McYN1gb27gx2uIvSDBmbzrnwI3d7lzDRD7
qQz0k/tdXX0iBKo19Nyjsf2Bk4Gpz8QKNokfExQeqQrclRBFqIcmdM0z9aRXlFAWgw2jo8bDyxcO
lb1b+0FchutFK7tDNDRuSMKRouYj4Sn3rwGRGdMWbNsc19VWQ4r4iM8mfWIOrG8Glqj68wBzd0Qn
rOCDPW8d73wfi3GfJzeUiudwz+MOaLLR8LazIaBdZZRMV+t4dCPuZf85VFZPScZY2g675eJkTGEh
YNS1XA5TiHkFCCVi9JJdGd7vyg5mZQomrdMEBc64MA50BzT+GRyiICDTHScoxeLGOUlj1GWVUfUC
dBJLIvjRq0Ks7vWs6047RyRaXifwxeF/VJtMy585TVMZPewvqMoUm6mpUMfKV22eMGzJt3vMpPKl
TvnbmN64BkfgdMd0x3WowmQWuIQAQumPYbP8nXIhMXcAgI46pMQG0O5Xae0jEbbNjIrUVwxS2kB2
/IdZe5uo9ahADD1cveMGBF55qNa52HGmIreGqdqrHFfINeRQpi/3FiAdh9U1ZMolJNZxRSXlah3z
3mVv80yRojebRbHAV68cHeQcIMQTioOk/T5oENh03Ee7adZo+gUUUjTTA91bkzKTV0JkuXrkBoIf
faisi+dGAjzXkWv+BXp1ceyfnI7gy86haHXTj5/H6cwzCcaATsM59/b9BhtbB4zSmx6tiOzQAros
t2eMyMn9dEufMDyWohXKn1NAjOuFu1qAYzSqsOmqVcFGGf/2pqlOZXcu++Rpe5FMW77A92tBmxvv
1GZmUoHnvPTqfH/M5ueFDL8gjJgIUK0Fe+vZmAl2xf2t9qrSH5PGrhff/XzV5PkoWG+IvpH9gpq3
/2l8WfZcsrk66iauSYUpkJy9n2BTG957Ojwe73vq4W3xVZNARbObyvldhix3ybojYU3C5tkHi05k
+ZGINiVy8Z0LXEhLMzrctmif2opFHW7v2JdZpuMMG2Vj6eVeoDlgD5iJDQLkhnn17bFybXeb8jfB
r8o0EdeRwW/qOPOrOFhqtuEcok/oxdK1h//BiEm+ggGCPAdWv1DHEol1xa9z781zOQHZdZqFX+6X
AmYzPMyWRF4xyca2KT85QLjI3GPwJjDnIcpCmML5NezHErUCT6q/Ax4hxA7pVV2We1IxPET05cmK
7HtQEB9iOfYBHEwV3YJ65oNrdUiJk+GxvHcXpMS8ZQ2WZkLaUlmzd7Ar1N/XvEI5Lt99jIV1kq4V
BoWpYz2VJuoqpCOp/DzIuULtU4aqcP+g24PX8tCHKDROiivJuLVTR26Efw6oaQAQq4IoGq00vs21
RhaZ/IzcBLZN12/kPamzNRwBsTT4vdHCuDU0IrOcrNP99Dp5lUnvr8G+Mf2YNHLpFplghelTLCRZ
l2a/d3S+mO7bJIv/MZlamB8XNiwder4iJJX0PpOCJmo77hWGA0aJ/KPk0ulP7Dbz+SpnYLo/CDSM
EE7SEx2yuqfp2kvE5VOfHatO1v+u3XTiwCSHQ65hvIeH+ZT0uEf2qCNdxTskzQ2PIHWzUBbSV1VN
RwSnW/AgOelvhxE++zz3W/egF5ZyI3JvNY5zp1Sj9p2BQumgZZDksyj7R8/ielOm2o6ART7ad995
stPGdnKQRlLO53d39MLJZrd1vTyRdI22SCJpig88Aw59EqrB3yY9ObycSgOhwSRemSOS1PNxY29f
nXjA4FpwaEWNy5JzteABzQmZ/f8SB/GqKK68zqMJfnFVvwOlcOEtAkNM5cQn0sd1DiFlYJwwfFOs
8XIHhQxZPEVe7X1fzbxf/a35y1Hy/v3fYZ8+q92ZWEA7rqXl4g0Y8wT4zPg2p2ge5Qcsq/CPl9R2
qeeIXhyWa8e1j3rtwCh4I72F8GknQKJXHn6gKWzkvo5qjS5a3WBApDsJc7D2zZ65VpwkrFi6qSLw
VcSYtpxbx+BdZwNRwB5d/gh/VmQ4qjVunTPg+9wUkxsUt1gh029e774u+JMxdU6pqDPLfOHtK8rY
MJ0R+h6tPRBTshTvvfr2ffcmQndVG6+SnCC9IjA96Ec6PJ+6P4zzK08FAALm4DMJY78n1U9fSR6T
QhfhHLqvGL4NoG/BrLM6pv+OEl4+bYbRt/R05O9p76vlaLl1qipanwuF/4HNXMGiRcOqrXtiv7CL
CCxaxkImc8YfQazRkNItAiWOPAYTpAj5eGlYUKjav82eiJ1/o7yFYROKJHKRDJfXhfNXmkAYiBY2
XmAqxta+TRSRZumVBtILaAUpE+bTbB4+NrAHkZ3Yd06KOlzw8BW+CLKbo/oeFZF5OW1/r2frah2d
R+qpd6h+BVqydPHpx2hR9kdwlPPoJZtI62O/kZyklRwL+Ez6QS8V4SmCU9X6u5G/zKNhzJenYYdR
WxGOOrIf5j2cf/pi3asQMZUV73o+9o8CiT2mhJ797eSTdrqfzHH3P+FM1fb0OEgkFAWv+m+0iXIf
qRvGXdyOo8u3HNLiGX6lvCyqXNp5A83C3Dl6cHIbemClpgRlwHdpw8xbzOBCyYlcDqMDqEbUEF9h
PI8RgwBx57zZvFtlvyQvnqIC3pRJ/9jrzdX0d9wy9Pj1K6gah8OmqQlgWn0n+2RKSEd8IDk9Fvvz
4OpNmllkN/dfW6zdsumj+2oigWDQhsmtAW3Z3FE9u5bTXMtQT0jB0/QIYsRGnGIbiVPbMHAikUGZ
JSGZN1YunCKPwLroc/8aIIu3IaPRJD6L9rFVcHxsDCaqh6lRri24E3CEv62MLlLE0qNjMf6WtqUK
bV51L7e8TudIwqbS5QHLwoSCQEdzepoHGefnlPoGwYa75C2tGAnGdT6i5l8C71Ux0X/S0NYcKAJB
s2Hj9o+RiyEI+r570nLzacWmZWtrAoO59N2QRXLF+7kc28MPbZIQVtHwSFEtj+re92s5clETJugo
IONsw3GyVyLgLLxq3ecDGvFj21BcNj9NQ29M5FJMEI5eSFaqxheOIm1JMOPOCPqud4V9jnq1J5kS
5ndSX4UjK4ZeEVl7ZzrFrAsSRsu6O8HwaBx33r/5p9JnbRul1ojAikUPnUgSVc7wtkHwXR6YJ279
rifcfthr7qGgideqGw7dIJ93DcfT8/KQbwj9VyAla0hIDZftiD5NBG9K+4uBNZ8Q1xMGNtetsEqC
kbBwDk993ku+gUcgsJ5zvCSKUXrJJEkE+tTa/wN5hu7HHipy3TJaR/7TSHFdLb/+DyYNOYKQjHXG
yeklS4OlqD8XqzkaXNhe1QFWaKPLHnS5uzYPchYoGG8L6r7pVYRA4yiebL+kEx26mTUyS1H15dpf
cdJNr4HqM8ndjRpPcpfnCKCaHQ79zaiOAelV8Bzv5cKOskOcF8zOPZbZnNscxXVT53EbecEN2zOw
MC8c+IJqhkUtMnqwxxi0htklVXfMab6GNu/z+szyiiVRtrSdWN3K040KJiIMG5pSFGP1+frjrWiG
hrT2FheYQfqy/yISgL/Kwy209mYLAYvuv61plIC3nY2T6TdzswPiMABymr/jO15F9L0aFy9b3949
CkW0g3pbSRMt9ya8jR+UOyTgW0RlLBeTuVtnuMe0ebJH6qfMshpyS5/vMaHirFyOmj2PGxnFykYq
BUavUgAubqLZkBRg7z2hTrmy3FS9zpKzYH6hnn+7fbw/jhbLXiiAEwvxEZ2qLgqyoXTk7NKxtzah
hsaR2JRiTQzRi0wviEIJWOa+2KgC3OK2rbqLCHD570jfDnI7AsdiIkSOF9wAoNP+3qAAipBEt6Tf
JfUCni2xufsdlwciraewvgxdLCIzGTWR1YIhLq4/zExWOmhetU3rZWz6oWfpDbUdM0gWiV4gTPpP
s2HMk33xjwHSffnFjMI9wDz9P5QMcJ4a8nUJHOecG50Z8L4n1cXQaumYricSbwt48NUse3b+Rg68
Kl7FmaY2JMG0LWzYZfBcg+tnGG9AJNBeTsh7TXpsA8puOjDw5iE6jWeBJ9uNOK5zAfqIiIysxAjC
8T2cfo0cVVbwPhGgH0r3l7R7xu97ypJXjV88NlXQGvEr5ujJ92qUdpMhuKj+jw/8BznSnBQzErkr
mxhAmGAxZoyfd6hxOA3fH8TBfYT9iG6qIKTg8EPp6dyZN1dzcWkSu0xNdfcwN023JGAYEcRfJpMw
7Zegmty+0DyqyBlKMYLAky/ujDf1CdHPmNN9DNvpSbDC8R9GH19qPjRwYDP+v99548+rLjPFBCVj
fQmfy/vaStV2E1HHJrd31OWC6ijqi6VeAgq0/75yGv2cMuFLdReNRLTkCwdQ0AegPKnfZ30thUby
ncKv9naqQdwpcE8nPrsesYxDuvEd2cmrfsxTSl0R+Sj4/a8Rv9oacmMOIKIcFFCxI1v2CEgiat2K
v3cM5px1jdrE34uCUqV3YRPhOL2JhlTB8UHgflwJZqtyBFGZuUTw1tT33ElezIoyuP2t4bcRZbH0
on1oonqKoGYaoK1lDNqyQz9diWqDkmrGKU15Md8dcIbg58DxOxDn8kQAYnnojKmE7oHGs2heHQLI
lXGMGVNJTfeT3AhCiSd2zAEPazCTOSOWRWbSZbFriwfMO8iGBgIaRHtz18/aT2wzp4zMjge4xEIO
cu3B2g2MBYzr3FoKT9402cXFLMltdG4ilSmC5w/Jnj791p4mhfvsM5rTyZAstlaMZvWdZVVAvjIr
S7j0RKObylIuH0M3Nheoj60vrRKD9VyhmmWpDxcP2DxXv9Ah0eu9ePREy7MaNoToFJDCK/86X/Yj
2+aNYeTlUrEdsADC+tUOIBupvmBzD6uubBTlTMToYTD7YEfXj/+EHj9m1O3J60+FRxeg5+jf2Dn8
iaQnvTcgd5q/atsxH+I0/cOKMEh5kgeWXhxmNfWp71weSX6pRVJUI2kDyI5d6CCLb3XSus9nXCIr
Ylowan8UNcJDE0iHtQ64xsryVpTjRGg5s4FjXrU5l/LcLnj1IHEhMmJb0BJmYUBrXPDrua05M1QD
cgBi5E7dGW7OClcEFsGuire5ihHKoDF7LM7/j4hKbE7/5YraSif/gcuwRWFwAmo1WOmTdPnE7vxL
6phP4CXgm6c7oJk/OmTGre+s2KdzBAgVVI5CvlAHCqilASt6hKJ5L3hPwqjyEbLKp7/PI+i8YM3h
mD1VfuAsbfpKHDCrFlgQ2vNrYMMddsFOyJbreqE3E8eBOOQbo8/KLL8o9zTznWR+sVoWfNGoQPVX
klRAM0mWFYhrK9o5KCiaFjrQd1owcaCvgILmSpM0u6L615lh9ahZBQepvglHTwA4uX0DKA9FpJV1
iQfRIZ54fpbL/shyza1Jw2ixR9iry15w78IGFB6VcxKiMPBTE0s68sMgxDwaiAcPI9k5oKSx0uGb
k7VajVfLKQTbnUufZm2XmDkjRFOmgOE6LbrrJPQqpMiqbn0XiL5rS4O2nvE4J7B5mgvXkyY64EPF
sqqdrbV3nuhFSBFmt2chi4MmvjhSZPw6CaHblypWdScDkBpfOLyovdYgwZPk6dqbrZb5dhln9Oz+
PfgbzM6Xw7FtxS8PrWQ87dluGOZN/hGNXSk05E7TA5nbf5B/nicKViKHPSA6NB1jEU3PJkK3hUoa
vNy57Kyq365pe/nToHwVpfawMsTNum2rEBe6du26s7zNV5lGyDe9R0/9h62eGBIxuk7uSMVs+mDR
0ER2G9PMXAq3+rNKi9QVmq+idcJppHFjt41q8+/ZrgH8L8E5Phg48qDbZNGO/e+zIW6FCO3H8xeO
SowflRWMCX1OMLOB2m7itryVAIKgNFWe+Pg9hpSYW5FjnkwcH69+Uq8HVWadTf2y8V4PzMPHRoMc
VqzbdEZ1q9sJ+R3yYRFAsqeA+d4+15gpCBah++0F3aOzLSL7X5gycODofj6cjH0rRT9B7OxAJ5Mh
tNvOEhA13+e1tYxuagn9Bar1Y8URlJ22SWq8KHyhuthV60mSl2QU90s5kgQt3R9wMX8wDak5Ri8U
DO/9L0zJIua24+GZm/B93LD2yc+jELU39inzrYESnNyU+yInryAIrzgMk3LYSRjSzEo7N5H3bAXP
i03wPPGiM8G81bXS5wykwI0HdFD6FcGOiOybXS4oewVqbUQW/G0NPu2uPs4HMZy1nA4meTvHvkpP
DGpuXpIbYImRU3w/QEe5Vy6O8eqrTxMXTmvsylndPuHLtKXL9Zu4/YMW1fZf6D/Iwl1w5OmWwOHM
ZbHNbUeazXfEaFActZ8B9Qdxa/n60xEWw27OXFP2OskRQdlT2lkbl2tHCvj6kaMJoubFNN7rYM2s
Ke894Te+hKPCP+BqO4rtCdtlZueBljCOf+B+dBsGhCerm89MSYoFs6fBSBix6gJBPcGnG9z9jzMe
9qmBnF2JIdlLIbHlfsuqfAnPJg8zWasVy4locyav5S8iO+M0ZzY0fhYc4t8NAeFoqIRHxA8l8rft
+gBzWUZmeO++mGw0xowRC/+AUqzChHhKR95VjrFUSRedrIugsRC8I6TrD7W5D0BZU0lESqDDw0We
ozmCHfnefSKcLmCUU/hh2DhnDFfxvbDxhcMUZgfdKnt4Ja+OyHYi7YAjDgwdjAjnZc3ZWyAOXVHj
2FK/2ukhP1EjTxHD9mvm+Dy0f8ijIikgZq3nY+e7xHI8lSa6GRjdJQgUUho4uKHaR4Tx3635Ahm6
hkP096DN1FOEPEuJo8stWE5B+dXRfD86kXn5LtExDLQVn40PZ0UxwjSWhVEINTBJb4QlYl33TyGu
84r63rO5rIFZhS2dAjolTlnmu3C+3foqHCaxB9giYLF+BgqtFDQzLolQ/3okV68a91yYO4oS7ymG
ycoKTXIpowwrDwL9kNVqrxBX5n6NcdUxMdhd/1bchISi5CwIHuZD3uf7dlPT6P7u/9bnkgxHs8in
6DtY6ATzjAj3dSsSGevLVA3SB2lt5fe1dZcQtFe6jsxDSe+TjXz8kBgeXTBg5TvEz1uLuofILmLw
bQQ7KoZ6i2L5ALIB8B0/qlGooEwNjaUQXcr3MI5L0M8DtJp+28dsCFz2tgAXxojB3ofkbdDMFqIH
yFsp/wpxACIc2WZ/XdNC6DrqxBtuYRPHjQh6KWq+DaIeu9lp5/XyBkQJGFCmYOs/aj/OUmNQaWc/
yUTZNahVBIBONk0dZfhBXpc1EO8CSs0SpNGK/9CTEcn2by8Xm23+BKyJY4wuqzC2WSlfb73mwLRP
IV6y8zPk7Ya2GfmiMr0r5kU92XiGNry9hZfT7qGrRFbGklmcOHOQ2V/mG5BkKSF1cQJ+e7IVDuyp
TfZq4we8DFkXj/dLbkCO+ovO71HGfpjo5Z+c2bv/NPbob536ZCoJqMFer95Xnh6D6h+7fjyOHmgG
6yXXun47myUI3cVtQgDoGSQvpzL8ekHLlQa1RLFcOpKCKWS9HYeKzQqG6GBjHk6BALwABbLwEvDh
0RAUfRyHCuIYtFtxsmVEvALmaNb1OZqwYRBXTZgm8A58kgbkvhPzx+Dek5pERFocw/it3BdcF1PU
FGywKvQ+CcmM/K9C3MEyydDfEDA9OoImNr19i0kEXZUAorLquNbFPlEQkOqqC1qv4M6Qb+Tu+bFx
VpP7Le4YpkSeDVQq4HQHIZowWgCZCGP+X3TfADV36SUlCwopuDhLjziFZKLXd6weDaY4fi9a4AEB
3R5s2ZOLQwbps0LE5aJObVfgI+OFwCjq+VlVJnO+QXsQPAziwyulj61DT+luNGQQwqezYk72OjbR
pgn7AZgFevdcpwKDkJ8GYIi1ZQXWoysCK76Ztu82MgtIXVIhtEaU9vjGMEjSHs48qBaRzpH72W5/
ZrPJaOVFISAQACTV8RuTv1hLhN9hKk8hDl6o5oqzorxK8NH4jsSw/q/3NNj2FWJ39nw9IuHXjTw3
pBmWOPzW8bAQ4isblvEWyRSXLEUPFTACla/ithuNs5LN6gk2+1Q0ed5+JVBK+bqeLz2/vScW2e+8
MxoIokSf1Q+j7n/0v8HekE02qdNtPWClvHu5i1tPWtKyLvNg4iWRnmPuv6aGGGh8bhGOSWOcZ4ov
JxSundFb4wWlWP/2Tg58LPmji+rD18+Aau/z/rxBAFITaXnu5lyDgX3IGWmjRwlcPgefjWnwQjvH
C0k/rKqBu2fbI3DPYMXMXGUFPnBUxj5k0EzXZaCBe0hI+vvbm75Xma91oVb+yeS0yT6G0agSGmDS
3w8zDEJzcQwK7iSgagivp9FGNwOXV96jkSQFGCFnNrBVZz5oZ+CB4HG65FvM+Fw9/0G874udKo8U
j9VidasBHwc9iv88B7XKjaDaX5xXFlTZN/6f+bJq19Pbk4KqBpWCT2fD1WK4srk1A4N19CZJhZXN
/JbICeom+qdCnxeNRQ9wAXHeLQBOJEtBpB/Fmy24KX51/sAo+A18SaoLXt9/yF2SXR+FNyF7Yiz8
zlbRTaJnmCWOnv5Jzge9MGYC09kgfXyzC0mTwHg5xTfaUDz7UXpN6r5/g0xGPhG1PjOMx/WSLsSx
ru9wvKV8kfIygxFQ5YfueBQWF9n4O+soVe/huUlmIn2wH4gER11pUbeBnHy2BX5sly+dEjgRgJiu
oZ1cbp6pz4J8QJMA/mwzu8/erctfWmhVDSfNJKsYLhwl+0Ael+2e9FM3ctcVjz1mswGdqT5IjP1p
FQKsj1SrArf0QHOO4JS6LvgeEaSejXBr7voeIN62urNUtlvV5A7YbKsLgOEHzjsU6Psc4wsLPdiu
WfbuuPIQoAsNP22ZHtNSwk2jKkYScmaAQbAPgKkCrqDCR6NHpbWr1q9ICj0EWHNIv96A7sKU9ZP8
6VMxla1GimMme/DfTt1aOmDqaOuWBcUM95y83XwIcG7gN0mku9K/+bAiH5gadiuK1O2H+27kkz97
jR5VUpzpCrAYqVXx92SGtS2ZjGJdEjA3JbFYksqj6/MeOjf3naNmHS5KenkwdReguq6ovYObBt2T
T850EYw9YwsBqE2qrN55x5xfAwSIJDujM1FKkIRtHbGgNsyR4SOseBhUXSXy8qoBZ5/vqPgf9Ebt
/mHczED1p2ZvVFR7kwoU48FTtGFEMlXpuFkSn2M3M3j0OnFQTUq7c2SIctatg1Fm4M59QyAZjHjT
BobE41SQgrzfXlytJvO5fXfNJOWz2758yj/THFh5LbWsEV5HeZhZZa65xDx0M+RG0sZfp7GZ3Z0l
VXIRW6wsdkUHCwt9N2Tm4VYWgHiMlt6L6f18nRbnvoDlJ5nzu0Xc3q9qAP7gfcJaj84JKiwsUvj9
1XKtxSJPyC9qV5ZHKWVuDszvGOaBeDT6nM4n1zV2U/Mvuy9eFFxijkgsYVjiU4VEdrqw5TJfDx7Q
CIVHeLm+KSey0hLMrlGs+Pp/bxZsZFkrMqKaBjaReCmER75atfWDxJCug5MYI+qXRRfaUbTfmMQG
71/kpZtTg8QULeaQbOTfvcRYpskLlmlp3PzMpBZS5lSe0BxhCMD0XkmtfPvBtK+n6cVQBMzboupw
tZjGU78BLWjWdShuR0iRY611Z/oAFKzXwc4Yeg2r4R1YalxEgupWqJtF+agigVKer10vY0LXOUPr
VIJCcy3MoJGps0+qSVliKJXCMBSDMi1liXTye2mJnjBS3YjM961WBeW48TGSdx39PNcuF+at2X1f
A+ElCAqomSo8lcXYvp5BsdUThD182tTgQwkKTek1uuMS8xeTPmjos2T4D7kXzZh2LiS8MVoBqmCN
ogH/z8TLx9dbKxtTH1LpwF0u6sXnUf+znqMFWOEOjEmwBHF/it7v0aTL2ogU+1FkN0KOg5QNgxsG
jWxiFwJ9hl2XFULEoiqrjCtptdT7RwS+DRqY9GLf68cct8bcMlGsWIaCTk1hbvVvkXeUCo3p9L5F
HbK3yg+HZhshGdJoy6NFr+k9oWnsmK6jdRheZLUV9Uvw+JFmOamivI+4tepqhUvyet83g6B6fai5
dgxjHqfBF5bhOhDrq00o+GaSjfOhj9DTaFf9k3xDxp82vMu4lCOIOCzeGhba1rHkg3BvQML7UUXC
206QYoHrcQa4YpvCPCwQGXo2fUz8/9UISMkD8i3fV7UZ44M9YtPiTTAtthW++WnvyGzkZO1YrCgB
Q/XjWeTZuR23Pj6SngtEDHJ3nTuGL5mUiNxpmu1Yz3+0SnB6GHhJU5a/0HGUHyMrPKOu8NA6IleI
O1wRRnf+KMkDPUH+jdE4cqx/9U/s+ucK3Yonnmh+UNjBjsbc/q3yStA8ZKWe9n7DOJk1iEexTSrZ
eIi/4z/veW5iknOSsapYYGedMisk3D7X51PLIBCdwP6SUIaSEBo1x/pqRj5Zgj+IZOVPmqCQWOdH
E7UmXaSNNNnw3+pVBk66m9wPB8hPpid4a2mtAJISBfdeI7HH2R02tT9CisNDQWDUWh2EL5XIaWdB
4X9sc1BF34ME4iXUPXY2MTT8PiTl9Ud+Fyzm875ObKt8igbKBK3IyiYkUbuah/Q2XgKm0cw36xhu
i4C72XyjS0Ofct72mYFXDZsFGHCUwwwOi4p0Y+8DLSCIb+XYtrGakrmHIzksMyXnmJeFeCRyxmCL
XUuc7ubZFCNMM8KN2suFARM77MteXkCV88G0EytTTukUBtZBOWMzina1RuMF32nArn++py8tLS1K
wvVcjNWZdxoW+Lqcfzg9Jy91TgBd0cMVPoLkgpWf8Zs9GO8cH40rMpsspQaLkuBo80WS/8j7Ltmh
dZ6y3QqVgnp0SNK1aK6tJDB7/Y8NwQR+Vw767NVL7rChb2JNlKYDZ65ysyEPqZDMOU5pjev2MK5D
n+zrq3Wrd3ApsVsjqTMfpgInsl2n4oLgbW98I1YtxohiIyL1jhCVzA+xFCwwaDfEo6LrHN+4Z4nt
Nlj7qPSQceEp9qpAWZAeg2ihdPIvH9S2P92+upH8Jnp2W4anAzJmLiFI6gInyTjMudx9D8M0oyAB
0NtV4+94+NAJ4bH4yxhnDEzENjEhAqWaOG/iQR06wN954MS/Ka+pu8ezv/J7zDSoBw+1DKLnDlX0
ELMzcNygU6F7SDcy6nqBTl9fTnHedVizj2udSaoq2h8cr9cTUuhMmbxKk8yFg0blxM5Mm0fDd4yH
0T2PM4/NGWsOKAAu+Df1w+Pt+wX/sE728yEaAD2mZ0hJVjwe+RtZXM+LJc8O60VCuS1g8Tw3mBeh
wvsRpM5knONoB+Fz2EBkj97fhaNFpad65NFWrwkBmFNb7/kKYEsy0XZ02xhyVSZpfqVjwnVQKal9
6WmDQQ2Os0qD8m5N5gw61bLKZaQmIdM+xifAJrOqgJLSLNeNHyePGS8n/CXOxZWGe5gFELiyYHer
nmgOdN/h6b6rB3w+IJfGTiGtf2bjC1YXHbGFlVyJCis2WYclW4suVk56u/VbXAZFkpblgmKL2/ss
cgHhejCc2LCgm/0ryEl2tbFyBzSfHlMgGa/rOl0qGi0/cFfZOozgbs9KWeZv89hbHsl3lqr5TsUE
pBBxxQU1JzKmhXouZbohAOv059b8zdVRAC91PMxzlAFcX8iJbxufGa6bgidpbhXp9EER2pMWL8ij
Hhr1cHx0qoS6/RzxHqHEn448/TUN/VUtECri5FbIkxr9HpHxz33NlshfWhcYW6k6qwMxKBg0jC5A
FBK8oYLnCg2BE6HmVmktVJIKrGWwdScgH+FKvhbbnkrnixidF2BgQB8RnNxWvAw6MwiPa8yImkrv
9/PQIKdUBpIhubviPqmDxGRFJdKY4puYJPuUVEmu8nGB8XOq66gG+Baq1OjUYU5F20prY6eWfCKk
qUNVMjASj11We7KMAJTmWT5H57vvIf8hbhvhBqxI4lQsQaXsGBIdpU06mOU4hfJk1PPw6KQb96Lc
ufSjyFmgXhwpOy5h40wF35sel3dRz+1ghxqU/d0OCtY01lMtX4hBuVIP3UgjgKEq+YEKf07xSmsw
t1AKx6+cUPCzwXTaOw4ZzjP5tB+qV1//QJIByY6xwWfUwg+CyVQvkL05pDx7KzcnbHBDj2oIrVLN
+wN4Sr52KNVGp8mnHHBsEQqbZEOHXZkewChzNJ1ZPtYTDT1hW0N+4pkVC7tR1Qk+k5enjsFpa2ni
zn7uAxGhXZ75npPfXDDu4+hlT2yza+ZSUV8Iaqx157CjWSbo8euCjjsYqcgfhk9J3LL0SOlj1a8h
Jrc0aTXlJrYQfZzlrnb4wvMzfYQg2p6VX6NUwtXPQMVxseTz6+2v4bFzpm9EMfPYhJWVi+ZUFCp1
4Gtz/+ZxAMrrJMDxuPezldkM6AO7kAtXf2dJK6BBeTSJdSCwiHtDoIC7cjVDvMrdmO6+XGVekuc4
SZCKDpApIpeFMs/Vhs5VHDDDHKFL2/D34d67iGOuHfP8R9oFEfFIqv/D/AFrnlW70DigqGy5EG80
N+vXW7OQgIPIFIx0HV0Bsbs6RxcEL3s7uMU7yxSJzu5y2oeh/cS+OLd6i5x0nNu/QbANs1a5oyTE
ifBqrLrQjdcg007KosifbUqa8rgSykoXrjZRjJ/bdo4sOJ6O++n4LY2wBFyFbAG7ldYsV1Svqd2s
TtDmY1nijtRFxplRQ+RO4M/AMiTYttStnIm92qkWPhniRBLg2qHQGFDaLSEiCtOnlxO9bQSy2Hw4
NQFB3EmfHM0k+PEbJ75ox1nln9r13SjNT5SjiHsfU0M7WsCLP0WIr3sMqQ6JSje63IZEYiGg9t7K
/Kl4Xjeyzs3vdhOK3N3MyLER8fG6L+AHrPTrGkbJq63ialoXEOqTTLzAUOKZkZifhwuSF15VIy0r
WliItJ34vox29rIiUZLj8x0cZKItlCO5yuFgtuRIQVEHwBTCSjTBfADE57ZlBHDwmvhsPu3alc7r
KNsWuVTBz1/2CNNPPq/4f2Zy2Xt7mNDKixabusJdVIYhrOS5cWjkpF0U0b5odg390Oz0ESeGlkqD
cdwfV2SJ/shRFT1h/tdq8V5bgPEpFwoXJuvc1rW01WT2C4CNsS+chsiHQytu8+i4LdpA/l0aX3bm
sF6uboohZZQneND2+3POtMLsVeor4009KGhx8XVj1MNwxaRHGMZImwNcZv4avKnVpOT9EOyxCZO0
AT8u/wGS9dNqSFskXzyzY3OdA31/hqQ26ITVvbV0CApZ6phHYpCuLFVGFaG74z0vHK12Z/tc4PG8
Zs/VANOFOTalz33fyK7tJqPfMaY6bYQSvLlfLAiaJg52lRhbutQnMAKweYkCL46uRPRPNodqhfv4
1HoAz268CNYna1XX2mojH/PDP3AkFptzVSgSigxXKdH7CkA5LIwJMmb6rrxJXekyJUVuMBn5Zbeo
RWOrqGDvrZ4yL+SyvqK2jBAcQKclRZmYjfcWNCHiof/Lg6J3jnKy6rHfe3N5zq3SCCqm6c1L4DQl
/EEPM4kO+I5Pjt9VoTnVE9Kbq2mfqFXMp9s8lN5u1kluWrlLcZ8d5wAtdLXT+HIhxu9QHMfyG40V
/nYTOghGsjxUAMcKzNtS2MY8WkA1abQhee/2RdjnkLekNvVvvhbbh4pxIhGbloT+hsZenU2aZ/PV
icXms3ytzwZwE7H6zVAwagfCXgtUoEYF9ZeIQt/QcZZlsICOCfvkJTJThuhriTuGmW+FCX1QLuJH
7n8YJxqQFMQQnmHqg2MDFWcb8vzPC/gZTSx24qi4OFZtNGp9LjjRo3wjWBdv5zGo5Aonap5g6E0o
pwl/ZZNxZPMsPKhCsmQPmlUUSFyMdKvd9RJVKXXQxADjCAd4dcXNlMTEzqk/4YuUddQYY54TEUjx
YLfXQsXTqUgKgjw2ZG/unV2eAtCW91dR9YvFwjFefRXLET1lt92uyd1KBzDWkbhMaPhnE/GHMtQj
4mDROdQPepC/waf0/2+ZVOTi3wnb7vYfAKclOhb2+XGR06gEWZ3/pz49Oqj2/GvM5/huU7vIEnKr
3IVx8cVvn2yDQZZJ0ZjqcmOMCBWyDeQ717w3dUuhYtKg4eyq/A3h5o675GlVmo0Zdyh20laOl4oo
vFocDphHW2jNggpy7Hn4krIpUdxkUu2JQE9Ly/Rfbn/bwKfG1HFpztD8FXWymhq69AfF0b1XpQNd
i94/ZsvRBj9FFO6FxfNYjFzcyf68s+mWg+CfwWi6BLSzjVy4vmp4/eGAcfc4qT58m5yW+Bgzq2JI
LnW+cA6NkpXmkocv9vYll+JdcttXg/o8ck/UkfAmQZNIooRRgb3Di/dBzxw1Oe1eFGrNgYfCAYek
vI0p/rj5YsjCId5+H0zCC7ldtfVKaDnrn+mBjMYJJiEcl3CBPPprd2EpBwIL9Y5YrhrIz76jV0Nz
uH6ljTM+Y85WWHC3ydPsf2jgEpeKRJt/vRkZhcGvadtOzrnF55p0vZr4CPnw8vcLCfeUuyGv2XJr
f0YAXa1+N8wOXNXGbttmkOmwBtD/O5Y+hUT4Fjn0PY7Qad3+asUq732KAf2si4GQdUe4XutZqtJK
NGTmH0O1SIhoaIKrLQ45SBTI4Dbrl4OsHA6r37uzl+aUyy4dV03b173n8YMXRXUV3WHkND+fiib5
gCaw3gIy61+exygwrXJr1O9jwsyz1LWubFuA8kmZYq+yI2XJ739dQXXBx8WSXU+9+L8dgKzN15e1
lrI8GRSxq8jpSpSkqfGpQlHLQbE3dzkEeRl5nUwktKJfDly5uPfd7cuWA3rvVZzsRliQv2Pv/t/Z
mgVwfAwVJC2Fjzky8GNpeBzn7f87A0HI2fALi0s8vZOrl+GAbDtZNvxO9PQDumScAEFtViU87dyp
bZDCj/tBLaiAsoMNuRvFrnvWqwU7X83Fkr4xMrtY4ikpQywxSoydCwS8IrRWAuDlmxJABswH6vxD
S6rZpHqc6BYrFo2PkBu75yQo7YOVWxZz2vzl8UfGc2hvSL0MfL+Ia5dfrthGeGkpcy+wxtMHx0Uu
YHqkOdyyIW8UnbtNkBFi63p5ijeIoQrKeNKFi54dutQtsJmzufDI7tNhQcE8SMVSKD3ev9600rp5
B+LtkyDgERmowXuu2BwvVHQ3AyJ4Ld0m6tMNKxqFnl9jCM9NKSJu0myTfLj7Bv9JCwbTL0AEEgdj
xFFF+9XYJaVWOVeKVrImOsDirhrMSqMXS7pGM/j0/nuAMS5yTlngF0aXli532PvkIApKrIKX4Hon
t2/3435IlPkjw+UY2V4unnQUdckZHezGaM+V7sqnHK3zhyXQDfJcSR5E1ZeCkOmfXNKmvkZYSa+y
L42VZE8OpFHaIQRmIzUenvxj4bxMgjqk/mhO9LxApqdVH1gUkdnHfqm503AKwkYN8D5ZZMGWoS7I
I3aYqMtz4oMp23wKfz96ffovVUJTl6b1xT3AeZdcRhUk3qJud2L0iCrnVeTU0fZ25w5MJ51xwmmc
nBdD9oBsWuuM4lqLph3fzAWfuA3/j7XBUpQPPIdZBSF2vi8SyEIJcGvK3Raj+8x8PICwlEGf/NnX
ebAt1YhXpsusp6XQM+lnE6kI9xikUKXYOir8E2vf83yhPAqfLalqN46lY9m2PxOV0iWYKtMak9Av
6USKDrvOVR2aZYqGWZRB8pnOJbCiuEYROW+pyyH/Tm6/JvdPDObIU1XIN+2LINKoQYf4JNeWzjgt
yGx0YOCn4tRQvoy5NNq3GfgYv/zU7KIHu1P+PbivUgps5yp4JS1uqbcX5unsWZNSusVlKS8Iqth2
/udn1RiKQDVonSSVcg3eAYkIk4VCL3DGlZdWrPf4MKPH6dIB3NAGIQ1Wu/w8qyWcFB8wxPuWuKj4
mvklmCIv7xNvJMA36vdKKD9iRue7Ui489fSHxKawJSyILEIhJgftFsCSl5+du+nwfAshsl7X2EGb
t1xmob/4mgN5/iqm+UMeRKYwsactTQclM7n9VFCPTrP0ioqbNIhDs+LbdSqH5FMlZFmDCa8iDDRV
qN2TiLDk6t79ohd7brgtcrcx/ntGwa5atdJIJO5poBKx87aAJFn+LMF/C5Tol9QMFOxXqS7cmmCt
NRee5vOUrLQ2IiV92RdmeLyKcm17C145NDeYaTSsPeJuIXv+y3vRv9lw17XEmcEMK/sA8S5oGG9r
W/dM56CjMakC6O04WMoAn4ECrAFh0BjPRDvxF0SxfyVOnlKTOWtoHI1d769g3OHh9H5JZfHRti+4
SOdYj9dy7UiLvoBq7OzVMdXp3LX0kxBwjU+HLULX8YLDaAoQyWCDvTqthQsO/yj6Gmr2Q1gU5ubf
AtvCcWzzV2800Ty0TUwmX3lnQaE6wwjK34ZjGUV++kiYaBBox8tBBfhDM9uy7FSOs3CiQWxMueBf
G/I/G1RsVXhl3JcpOB5A3NaePzXgYSR2nOD8HHuvhWt/MDv1gmifeg2f9kxqFmab8YzUaMXD5RVS
Ybs4P+naTcJxa5juqdNbKo0ZGbJAPenK2mFS+qhyv51KeUHHqRXsAlOEx030DCYdn5Z3jXCUajtq
aHxpQ+OFo7mPmKfn/6UdohrKcE+L53DN1oMMaYlkXyrtxKE5BAXul4B79ZQrnTLt4S3SgUHbHRYj
lLtSs+m0DydfZk+gouEfYFSJsp5nHfCN9GI57Xltxf+l2I2DgqpRqGHwWbj8jmXnmoJhGkfIk+R/
4LgWHVYoN97TrsTeV2YrhlTjNskduvC1C7/XPDoi6g+jSXbscvnA6ezOxo91i0ArxoryqITnFU0+
Sff9cSK5AYoW/jfGKGn/Fd+ZX6pNNFgNc6/c5kFoXkgP+/uOYxQEPtGoxTt8vXbscHtto3TR6bn8
ejPVWQOojmW0NYgIf6DUSkQ2dpRS+lEAmxpS8J17crtqan7wDk0q06yu2Bp5IzQAb1CBuZiN2C7X
juNvSAB5Totq2b6eo7Psl0JGl3bnzC/HH1s2Ms77emmT+tMznI1lY1m05sS042YCzVtwNo8/ukbp
UrL5DpwQ2n2Vm+lacAYVknndtvbjb4J0ePfZP2vrQ+7O1DD1zgssRlJf3Na5LtKOAcxIL7qNVAZ8
TmzTR4kBKLYmUln5gSL3DzXL4iv1q9MjmyzluIHNQx3oXhRupA8fztGWk0Zuw7rLggtbFNaTDFIN
Me/VH319WQx5+Y0r9MP9urbw/aF6HpN6xO5GCYLI4lpav8YngpmTf+6AqWyOKOUgDEZprUfiKOPs
mzzdRMMBcSxy75hh5IB5L89RRBgD91OaO4D55K8CKNmdln6I5ADz/9bAS/f76wrYXkiBv0UtDwav
NPFOtUwvgn5C1mxnIgtiSw1xujs/yqoZk3APtidSpoGkexZpOqtURncbA5CRJXu3+PC8PprMzeyt
guiijJRsb4E21K95G4vmvKJ0O8Vj0NpP48rJSkh8jmrgnsAtxqBDwASRKhl1X2Bntd1x6MjEQVd3
wp8jRIne5TnUEoKTCekxn01wCaSyK6G7ap4XUyJgFxbTmcVIMA+Xu3zJYyn8g0ZBBPxrp8orEhzb
iAaXYtRTMSfKwbMSkLPVJZXbaJVCeQdvyRmpm9vjav9nwic96WeEy/hpS9aUxp9TF1dv1LNtBhkE
ctk2WvRChXl8475vy75Wpi9XaRfKVV0LS/km7HAAL0MSTWdbHiAppg7WoUxcQYQSS8oqauCw2AsG
csXuMzD78CndkfPHnM8z8MospCPY3KGaAWmF6ZtzecLFYuS/K7+prr/jrgq8HmPZDrnYjDjhAMG1
N/rw6mGx6UFspl2YGVv/vK38NzowlC9iFy0D50NtYz7M44WqmeE4d2D4oz7+sdPOozaY87JPJDwP
wIxgfgjIbXRZBoNJj2bYz0XbIs88SNfbnjaRbVKR7DmyD3AaBKkSNb5HQ4RkVD+a+U3JvYc5xkJz
frr8yopywM+g69gAXswZfGU7dA/RZEnZ4DcCVkAzxwc8beyQ4AkVfcsVyfNS/Dslk1jiPS41kOQ+
mZ07TyIEWQ5Mz6w0dff+I+oI06ZMxdMITBoWII/H2w2EEfrq+TowDs+sxtpZWecB9Suh/6CApy1j
uTRGks7XEJboUgtKQeWNtP4RuAI0NKnysE/RRLbfOF2NhyUi6VuBw4jPj5KGWG3IGGcOpVsdDOOT
+yXQQyal9lrAkL0aU3oHhBT3WmcOocFu5dT0FEvDxVc5n5YLy1DxsHszGI/IfjzojXxQJHZ2kjFK
finmKEuFHUJcAyb+wLsrjSP+dJyS5FGbBAjLWgWgYLbBSDxXn+Iv1NyK/t+rBepKJJEYtlhkLUYl
10j1tbAJa6+4R+1KYL0Vue4YGr1tv1cSnV4u+QWMIQTnCZkM5+E996IlBllome1hv30PYMRGubD2
yBpcfV6W10+TjL8PKYV9UDSuxGG7q+eTRjl6OSWGWHW0WDByfCWZFkzMtBJtd9S10mVomM67vPzp
ZBJcaxqosBt8Yc5MedpirQi8yUE/lwP3Cum+mpACL5+UDWuikJhj950A/uLipSbp9aXRWq4K2M7P
oCxuDEe+NtMGKlTLDl/amhvbglmoQfBcPgka8uTX7kQ2uHtca/f/uSFhR43GGqq9Fz/XskFIOF4J
760ncepEFwkbWq2f+650FBKr+nKSm2Che3W4tp0oWOWLxnBBdOW/ptM2tQNxR49l7Oci2Wm7NS8k
28dbwJfQZXNlqYTKoYJDuqwVj1t0doeJe7OUoMinSMAVF2dl/z+RfD9I5QC2UYLOfoR58Xmk5kwC
WhPV5wC299P0rzTqRJuAbFjTDRLosnR16aJV2SItWzmfADV+Ck0TrWEHVAvwklkhsoRQ6cz3+AXu
RHrTEfabis3iQkU1sBL09R2vRGsEl4pRZZWRdQtByc6whm7JNg4e1msdw3XuKN8EsJ9DtJSiyG7C
Fk1DMJhdjYbekcvP2t4WQZUiNe6zMBQj5p2KujFE8pxdyU/APwbSucTMePKZxA5sDTYCJaiqX/L+
0CSsb9YmXkeA8lXYOE1Nzos+AgZxcU6hqxHp9cJJF5+onVzXBWCzt/qys2gsatpQvwuOLbFIh4K8
dAyJOn5McrW71sfAhcVrpitlxESKZ6o7WR6Jme6/x4Z1cgWKtAJfKEFtVsQRjj5/HuG4OUy1nsOo
tfaptYEr8uGJ+yt9l110ZuCnPwxX+k7G/Cxb6f9wzsMuvlBw9WcUfNRotHd/4BP13m7ZgfXJJi8z
nGl/W/2qZdba7Axouj1XgLvNWQtfKKJscd+odn9wesxVCdlhgzOUE3Nw+lJJDYN1eRNp2Db7N8NM
SCsfFTBrye/R88HO/BBjEFTlV7/NWbL9fQfBjka2D8gSqJiJI+bjNO3iIJK3Qx/vyFQiCnkgZcA/
3HHP/dcaWe5MdQaPl2DzPTEZYlBdKXfK6aZBlQeH9v/MxAd59k3yNkU+XP9e3y3jQAL7/h92URoT
A8QikEdxcGgh5zwvo8X2XOB8pZv1rqQdquzh9EcFFyqtclQDVggyHP1Ye/gPVVW1WHR70pTtIHzK
7QR2HOb0HTu5U63SzGxkGxavGi8Rf11la0O4Nabg03bgz1F7hwjQP6YHeWCaCt1Ugt/y6SUBM9L2
BVVqEQ7eU02xnOr62ECNyDzsNxnHJkqRGl3IP6NhzTF4vUKgqCrB5QoqDeO6yICteUCJTteXWwWy
xP+ormhMrigkZB7F2/eb2psH5Bntq9FADjTEEZtQcKx7OYLSG2qKOnj85snYTNeMtFZs4/rDX7JV
KCqkOnKTtLolJsakbjVz1Q4Z8hsYwh7RD/toS5y+1ChHO4828Dc4gEwZw7bf/dn+V8LY4PKVL6f3
/+c3WtrWwgww/6QXsBhtaWS7H54UovK9DFNEVc0JEhWtd45J0kLXE4kn9nyQdM9N1M4pLrxtj8sI
ltj3yCgDgEIvZapc3Yuv52qP7ZvSktVKUOG/5gBygUaRVQZm5NNKSkAXus6j3jOJveTks1mfMDUi
Gbh3NhdZ8e3vHNtVWFnNO7GhiNuO2xvO7cmuKQqUJ8W7pFFSHMKxn3Rvl8/MHrWZr/Pos7CrJMKp
SbfW3uA5fcFhzu72a0GwRg/+cZA8rMXZyAQJ1bsIOImnJ1JsmfdjihcEGolb2/g87TPZbZp5yn2v
snIafTvagP3AuptSDecUrnJoevpDaoVMponJC/87AbaM+PbMCRes+OEG3jVZWz2ah4TFJPpbV+/M
QqiD43Ng5MXVTCrY8Y7WIEsKlk6MxSmiT90CmzYk4rgK+uSWm9joAMuoPwDMGY+Yjs3mnlxKiI7G
WYwpfUL/qPrDT6RusikK1aN/qYl0jXEqulM4pZo/kNMErZ78vwuemeZooP6pqUfT4MbV2X2BytER
Yfb/njPc62cZUYJQh/LY5/7WlemEwonCkJ+AAH3ap7cQEwpO3rCsA0/PqArHSqWzfuGbllv3sltz
LDDIPJUBbai4PJA/mX5hBTR2Ur+z/CUk/LnzgldY2y/BGLwkYBOSe6rtgYJZ2yOIzG3FXd/RFWwm
SWl7uRLWi3MyP6A2TB4yX3H0r2IO+9HRmRkfdXTY3MiqWFv7Ic81/+tADmz0FsKvWdPoIj2xQbqC
q4GYDH56T3TShnqutBNwkHmiDfUCTKI0kSbc+kWkYLsc12vZzhW2QhTpXRpKK1LmZaTYjp4/uA9J
ZNOUR8Pif0byqql3DCxlwCS8U+A/Br1nIOrjaXx6fSHbY/pycCERBh51r5kxEG2XxIubwpZlUaKD
HybyrRg8FvqzFc7LsO2WcBOMAziLpW6dNPZl/PCxI+hmrFNOk4cb6Xx+hHhpNVrXkktZnB9vsDDz
Hc5pNP6gKdvSkLDptZ6tVD5NZ/cqoMK6iOuICckeBd/KhyZRywaR+Z9Qp0c0eapvGACoszBfiWRz
kZl6968fNtCgd+CjPt23wt6r2di3Az+YEn0vCYDun+w0ADbSpqJVkvtZvE7W+jhwr8I4EgLbX0XO
el0wlN7Vv7/sfu7JuurX1agHhdWwjWmT2dnYTBkuGANwtFc8mF4GVWvJXFT8EahwuBrriGHMbPK9
Or1SZgQuoodobevYLpkrUruSpbVaTD5QrtMzFzPXalm7HPNB8V0mJ0ivAL8sLMdn+ZszQwN4e631
Ij8ySywR+OdmXRpnO+rZuvWXEgPiZhMv8273ZsBMuuAEZZ6YhwpwYW+awD/XyjTrqRXt5+KwrMW5
QjZzrz5Vu9FHxUaU70TyZMKJjCAbYdsU76mbocP8uFTNXDy/NG9WKtq/IsgMbsBPlXDZCZl7fTUX
hv8WB1k94T0FUkXQzHmXFJKVJEGrjbPzVXD38fNmM565LWNaUwxfAaG8DPr8pZPgGcGZJZrL0F3d
rcR4cFDpCSNMu2eMPYeASJ8xPMtArHPQ7Q+spEnJ5OPCaQ0nVgvF5mS+y1N+JeJ+ZbLFFiP+1Ckq
KwOTSJy8XWEKj0YyAJ27vfTSoNseasM/qF8F7VjOXl8PSxcFzsWGK+CYIBnPs7PJLJIycbpy3fPA
yf6x9AfVxWcjumjWRqZj+SsQKoqsn3KsNz0g6a2kicpbf/HgJ1ywizouGJtr3EIIgIEPrPXKwZvw
Ojz3yW3x924a4yJXtwH6lJezBzTbvqPYGI1OPG0ccYYOjt6h29C79GIsAW9D3neutedtOurCjbJf
Lv0blzb9ippiL3EUrch9GG1cn0Z1DHoPbgoHazwjJMQOYYokdsbpd975ev11ZNVBc+yRqc2Ixk8n
+UJ9lxzWImVb1qoG/QvPTU+0PSK6KRWg7PhXvOQJmEKbQK42qzOQkSUZLSZf1Lkz3joPpySOSqyY
Oydmi70gaMPyDLu11gAm8F6SlZ6QoHe+oFiDlJysJQYv3VMD4eFtbYmhjcNUN41FFYOkc52Hz6HJ
qiV7cAl6DB+LahZ81kac8O00iwjKbMu2LptFFOFQa+l0hzvljd9StedQjGUtjXx+2Zvi/3KprlV2
o5h3+e+byLSJj9oQ16BGcLvFjsTAA8EyW2FhIZT32jU2rPlPL5XOoRSNEFCCmAdMIjyKer6OOUUk
8ZCt/SA4D03iphIx3EJwzMyhlja7b1/CIrU4vyDXZMsMCmrZf8nDPadpfBTEZdTIKEp51uOT8Bn6
CABBVgBrIkxC5c1hoaOlb3JqQODv5jx60ZaPNCQ/7C0wrRlmPf2pDxQt7bjhTR8kPfzG//wIX+x6
X605unz7XvXmY433m0VkKqxhlsWcpdEpP6hDpSl1z++2/Px5TbFk8t4btr/vrAZGstE896sw2EJt
KWV9p2lEdxbjTvp8FOGKyzpFrLe9KVrdByN0Cj/aFCzB0Ecgvp90ZmPZyEN2IHZrDkp9uS+R8lKb
CeDstaI9lv9Cnz3w/IGT2PlAE4RPl0oDyf/6aZTd6F2WSk3Thh50QbKP8RI1nKg0A2zZZ3ua+C25
x/utUeK25zXZtnDiB7HQAy2qYbNddN/DOfb4BN7+NLEfP6vbrczj0YJiy6GEfXJWWIxJl8PyrHFS
SacgjzS2tbO1XFl5TiKkM+belkr9iFSbEf/QMdaEbRFuSKXC/SEgoj1wQJ/yMMDmlXu2g5mJnz2Y
mLGp+bKUk4HK/SUdBoscmTnuBLwyOpNL9Z1nNxN1A+XxP2Zz2+0DImheTguI/kKkE+iQErlbHRwj
+MZ4CB6lmyhxEftFBMxkRUpmjtXW+Y+uDsSliIhEPb6KK23UaZXvXAXBeNrdAXdVmDzYuzVZYCYy
RytelNmA2ceNuAC2M5P0KfPIkzf3lGD63MODxNmpfJFKB9V4SrNDn7iTgXo2N0/2+LDSpAkeIq0D
H6oixGT//5u+vmHN5IUHfwL6QxDyDPNYWfjtGDnXxJTlJc4TcIfz9W9ESaFZCxZw7wqnhYWhcJRr
W9AarAOfgBIAcLDbcjYzoJaUf7hPlWM++VKJh29jLT0ITZ6vTHAB9fUbnSofiGbaEaRrH/0vyP/v
0FVdTkOJKHf+BTyFbCb2cFHTcXsXGtaVkUCnFxuVUsylx4hhpMx1VhnE/lfweDtc3pnCdKdYu2ai
u5LICBqyjTtKF1YQM+dM/UTV7wkcr1fd5ZhLQSxsQxvoRv/psXdE/d3ty8MjzeLTVvjSzuS03iqP
VDxveqgi6ys0BhfADo+J79nQB+5rKpwqNnagf0XtMuJGScOFbBAeKsAHLrZLlCC5PWBbUdjNkP4K
TLnULjV1aHMpO/fSSc0BYfjV/Bi3FDo2LW1O8qWplMUI5tMMiKor3HoFBIJYcaCgjI30QOIJTdqB
ULIS+x5b8ldh9bLmB7UAV2xI+Y6MqvMcYPIieoEyaFAIiZr5Wg0p5RbGzX/6h6/Dx6Y2e+CjoyO0
Q+6fnKSyL/Rfrzo2W42ZyBw2gSBjqq5fmBWLUSgT6irnvNzSvWsQW6F7WmjaH28X5lKISBdsbhEs
pjyrZPPxeQZKPElEB8Cq7tkmGtlp2Y6aIT4Oa1K2cH6tuL6ctxR9OjIbZPxduuzvIqM+bkPq2B5z
fQFvxQ6XHWxV8mcQud1P6mQjjZYifjfjBVl0gREW2pOIT5dwS+j+3P6J5TsSsixGNPJ4nqnK7j2E
tXxqVzl7m7VoXBL0E/+fNdVdBuKAzCMwwVYzk8WqzsE3wMn2KUvdhSJ+FAbpIoOQa2CIPWMZv/kf
bJVeJhfiOhuL1ncJNmW4z5nk75HDijKfHwI174Zx/1Kc5NlQh9rAXLvreOikT/bzcdm7Ud6kZIJm
itukJhw5wRH45/2RV849Kl5fAu8sVGoxYSqxKC70udl15FzPPVAjWYGekYD/HfQFD1feSUKwZ80o
x8aqa3sZmSGPSJw6WEbl+3xJb75z0Z6cCi8oXc5IvkSiDTTQ+g6MyT+NiuReMN75Z9Ca5s6lMyke
RBNlrVHXiWgolNzuFp//z5sU8B8vrFvqyy57a3HaKdbAiacTlsipCOhDgat2W6I5Zl8ix/1SqEd8
QfF+nsndi45mJP1ZYQVt4wM1MoBeFas/ty3R9QTR9uDNEn0SgtRgUQXcWWe8oNFAIGaaFqaIqDv1
wIHhWuPf1g7majFKfkMqViFQRB9ZO4sVYmbaxvyI7ZB2wEET6DaA2mH9+Y1u9tim8oiA8n1DAXoG
nXxZMZQ8PpgFJTb2T3oTIdUGqnbCQji40/T/FTNAmDO/OZDPsZik2xMArXq/xlvZ+A1GU6LL7CSr
S6f64sFljOWiEfhwnEzr2AIQUWMQxCaLtj3NQrOEdYXPQN84ipz5pJ5ta8cXUnHkb8p0RWQ2JO3H
BICbX31Z+5B0ws+IyRL+fF9EP6w06VKQDU2p37F7AOjA9PRrPiSPYz/xE/rmAdIxEJbKWpWH+zeq
K9WdTSqW517D7JtOY7VJdn0qdkw7kGaUIfjJ01FUZp9czyZkFjS7IGPsR9FJb9ebGNPy466KpFAW
Psjp4V32JXkqzIZZLWVYcXkWxg6B1jUe/5s2Fg6NeANrRcUFDSGqnKG+wRxZX6dzba8OnWRu4In7
6Q7/j9ngjcP02JhZ6WB4ksdiXjm4HI+4XJwcqsz+Gk8ocAXBQSg/mnDIIyCczu0FKFIdy2zb55xZ
Upgkz5BUseLx6jvIAowUCCzx64cJI0esOMn3RQz9r7F26SOXV6Gkcb2+eP+vAlnCFGoB8t827cbR
EaiSBs5unAM2tzQX1/L43DD/HCnA2Y7n8opEjq4q/3gblCBkybu6KKHmF6sCmnhve65EWJBbymrs
uGRTO3y6o1K2X0VGmNCnF0lANvWuJsB0s0Rt6fpPvmiSqkMPFvRgT/HliSUsdaOEkOrE6BKMRHzB
o8Zf6Cf9bVBhrwex2N/5NxUEJpWoFxlIVhtfbO+l3Z2f74eozeLqjDSZ9oWw614ac/uJFcP/adB3
4WYCBvZJEVIpyqgcKqgyWK74preigDvwgdUNJCjIPemOQ3TK125je+EsGkaEHiCKOAWlgOqyBVme
acYDe2WOKfvS9Z3LUL7Kk/8A2A80/sqL5/X6lqq0OpNdwXqoeK/u9yEvVzsjl9yIkI8v0uhNO1Ad
kWWUsuE0xXLNKiiGPJMsIoy5PeqThF2jhqLxIgHlj0wtcTzUUVSF2z3Zh+cTCeM1JARjEyyqHC2o
QbnAznch9fUnrGa0IpCETzMazjFejV4wBYfu0SDRx93BfAohsXccPqKoTmOJHy9qAtmQWRL5xPDp
P4OseWx6DOQAPOzgE5KTqUPbG+knYBQVlXg++67A0eQ53PojfR7wwU83Di65XLhI+Kf4+ARQYWyY
iqu8pMIITn9ZVf0ZjeB7NnwlykQyGM21yEX2tdlsN6NgNN3k2yzycjYxrR8aUbsIwEol6oi1vMlE
uLUbA0vtM9s8XSOsUxyXezEP8+NshWB1Pv1gaPinEVoY18TvFBuajYjpnHkQgIq9LULNJfA7vkHU
2CplB51NJHWnlV59FigSWHZL2/IRBMwarnmdDLLO2kYvmiBNpRD2NIq2A6YQiXXSjfBj9/T3FpJs
srhDUEQnIH/8FhIl+8aR7yXi+mGreP7a2CGWIis1g6tI/vyEVZf3v2OPbZmhmosvrokQTbaiZIdk
XiuhDwLhiLrvWgoV4H4jEihCVu2y46gONHCbEP4m268XdiQ+vKd65xWwxo6gvBLv7jH5V62nwI5B
FL3+F4I57axHGrjXoFoO5Vcztgmw5gTVyfdmnKiy9cNYYk5DnvyrDdhuofFu9TExBeSJ3BUPvg/e
bM7j76KJRVLnCX/gjjKP7kQ8fVZUdD4X0Wr3KhWhYrGkwQGSNQ7u1MWc4+4LtZcYF6tuU0AcqFBn
Qkmk/GDvN+KIOv/4XAMQsjrl805BclO1Y6Q6tMmIFIbz1v8vmAxm2dDtuYCDfPn4jWbitoK3EDVA
wZG5fTpn3jvyUcoPQNrInc3S1bJonxDAcx3YFrjYhOXgEu+GGQb3hCw+Kmzytk/iEwzhSi9zNG01
zOU7jVuxUNKuExE+b87LioPTGf9CEeH9X/tqVwP6eYO9VGM0KJ8YcGU0RpJivnzoTwvO1kfbiNZX
CdeEiYtsqLft15NQR/l1m7jaaRDCvvApjdQYafM3H5Z/P/dZOyc1ajSOt+uP7j+ti5jyH1GrgQ18
JsR2uLWvfhSHQ1wvYtKm1Rs5iXZk5imcDKxDVX/O0IsvWS1M6YXov2SwzuKueZodAsxeOFWUwN5Z
lnx16vnSGneXpSJl8vIeckfT8wBRyUVWdqLNGyh505syGe2YnsBYdezCjHRhDaIN8oZs4zwzoukq
S4aZO50Sd/tIrt9wbDSNdPRWiE3nHERbqYcGzOnNX35Aln253KzKMXWnBFrLA1oAK01mIU9SYWPL
s1n1GN1wiPgKdY5x0tn9R/Can7+9FIOKNdcb6OL/PrMRRFTcCRJz3737MgtwtjtggSkoGnWA53f2
6noMk/L/lN02VABl5z6TzyUnZB47yak8URsHwGJ4b4AG/uRaOf46VIHFRRSBA8lCaRs/fMuvBrQA
QqhpMAwOt+T2GDSWhTBfB7+xfNSAz4G3S8ZX9lAoYPE9UafgyuPnXbmRyHv03EBhxwbI52fVWT0k
PyoMC0YDHAUupQCUHxyqCIWgoFeUgFkgBy0VthlzikYMn8MZxUwoVj08bejas1eP3CC0VnFLKvDh
YfuJXJg1gQaL+L6nVGyM/ksuIll/00lrPw9Fhv8QCrcMMeNtpeP6ssK2oNufYtP8ZrDNY0xkOQtK
h6Z1IHxKNJALx6qn6ueEVy1Y1rEhlYuLGZ3glWxwH6tJGS2DGHfjzT1LwOReFlUHyCrLN1dof3SM
NMDEr7H9EwyweELqEZVYllSIDa1k5Tq6UQNw70umrUgjwuyXPWM7WfsrEA+NOQrn49yV8IsbuBUm
AHBO5Hf+H0FsxLZZ0hU77Mw81u7nRpSSdbJckci4UG+fWvqXU0JC8UIikuIuTzBZ8ThfHyH1g6KW
aAR4YDq+OQCZOShTjgbMzm+YK+xvMqD3dHqF6ShpRWzaBtDxl1il00SHh41jmB9qfw28IOtlW6cy
czuK+agvbQPhIKH+zH8tWJzOlIvGkBWZo3ICVSvCh4RVdkrzDy5PHGwqHT6UWgjcCo8Dd9JDIsMZ
IRY0kCgf255yU3dPz80ePf+DvSK5GE8IIHOt3BmO6VX+EJYCT4763J73+pQgbhVOTf4jxiVTvsmG
HGo5pUbjW8dXmdnHPrDMgO57nPH1WWKu/KvEsd/pz7Jg9iddp5HXPb0aHnzC3MzxLzBzlD3d3vx0
KLT4XfduWMEILjVKl5qdhr54uEPLSk08HJiAm+csIQ9H/iofLGS7ISUH6tGk9/eolS6RxNz7n0nP
MQOOIAMOLH9Dj3eOHTnokcyW9LKXty7nkUe42LVBIhVO1I2H0UvxUnEb6YsCfI5MTjiWOo7fXKuV
QOudA/fKq6fEpcZ88rgx/TdyJew+v03JYO7egmUPyT9kOw+yHVuROJDrTDPNuf3LsCgeX1uOYwbf
xzBxpqsCd3oMehaGhW9EvKKLwia4iF09d9ixi50Rh7yDi6Lmf67OC797NdZx0a47YeKNVTl6NPfi
WH1KV/ufD9zOUoy8nOIkfsRJvb43lVXKA55zI5s8icehK+fClObtAEfWYgULUdP4mSLa0+L1GVAo
SmB9Qkq3/K+irdQPJyq+8IoO1dc9Oez/sAEBf0SeO8QYPrnls+EMC6TeEBtggDt0oqd4qQqe3S7r
A4xkVeAtIm7IoRPkRmUrumpQeyVDRghcf08Ku6VdJ2+ggxtTl/JsL8RYUTkpWvk/Y4v5HKLD4+7O
FZEgvdzfn/7c+9uHUVWgJ4eLAA9NgRQHMLkPuIUteImAeurr+SQhyFrJpjo6MYDRgqMDI+xyuzXP
1u8wiKa7xLHmUkf2REF8JWi0l6LGjU+oUJmg5eWQCyZ/LuNpTWeZYeNer1TJfqwcK34AErceM3gH
vBTqV4Le/Gl+MwSS7MHdPT8rM+2rQ1uYGS8S5x6ipMkgYIn4AmosFde2xvwPEQoXIf5bBcwflyFM
6q9UNajVRQ+6nVAAoqhFR269R8DK4Ko9WrPw8rruYtTsFhyqur9XBQttbjOUqysvVm+0BbDquVEI
D8dDN8+2yG4kH6EfVl54olOSwqkgmw4iNiOwOYsQZ7JlM/q6Raf1j4bMPTFkyguW1Dl7wA5oWata
zVRmcKqnJitU+BRMvbFCiLmHDVc7NfEj2y22tjZLAUvgknOTGrQ92jITmkeKHrzZM7OhUrFUH6oN
mNwfys6U/iOt8xDeTrwLoFCttGbwBruIHBIUHSHJHqb6kE0h3RMvo+DWACmN1B5m3M7sgdIs4QFn
lM1D34VoX3nMBtKtAUFRdrf841YJURVdkSLH9JbTLn6IDVGbgbIHwgaBs6o7tb1uL40u4aoNCbGU
QPy2GKnQdzink/P2AZLzbVExJWIBN+cNbx6tL0wLWTt9c5eWJRfkvE53BHRKqXRpMuDzMeORMW+V
euTLymeeKfT4Gv2kvyvTv4e23duy1lIWoR660ZouEjhmHajHWjVCDU25z7Zetsa5plro6BIRSXob
vjPvnc8R6KK7SMtsBW2hIoaKPaiJmObjyEhuh0UnVWjgjn/r5V0b1sPTSwKyZ3B5vKO0TQAX2zzc
ElMsxX3W1/zLhBe/6BxLMgSOyDqR2VLdr8fB7H/KJe95GT7NwIVTy6PF91RzaMqzER1A2r+dKqVb
x2Q6IZ84Txx2p1C6YbdhNQs1J3i9IOiylaKk7RF/6v76ZQakQwpBa1DXrcOKn1SS/Q/l+Ngei0bC
Qys36eE6fTqy+K5QEHj2MHMWEo3ng/jwV6ohAoO4S/TExhz1xqcjZOt6XSIPrOhecUUvRiMJ9dnb
Ug5tvN7xhof4Y2k4yAPAHMcnKNKiIlyJRPbTZsNtCwRyB50YqJiRckq/WaUilVA69+yjBO+k0h11
ifBEHQlcsndW9sgfA4EhrfG41dL7JZrxeQaAoiTP95JxZKlxukSdo8DG5DF50yXKVL2t5gnEH4PO
t3wNKf2PZ5kpzUic3ZAI09WHx7AnZ8RfwY8z6cffwYEW2l1angiw54fKWd+xOzm7Ciu0p4V7mCZr
28bx/P+zBAz2/b+qDT3+5oBDFae4iOkz+22phsDDbaRWbhQzJdcFl4Lsh58nrRX5B4WTiuP2gGmu
W2wAR42YJkJQWIfuaXhdmowPKC/mhrS7lZMSsb+sEwvEyFuIFrQdcELlo0HiuVj5UudlDEcJYjXB
FO7dwNKU3ocRfWtjj8OJ6+YFNtAtdIZ+KxYP/Vn2c8Z2M9jbKyReCjK1vmkHTnXuRr1yV6w9+S4S
gbNTk0Qdy1gRfKCJZhxtdrJPxOYVEJPuaM2BFv7KSMaVxza2p8vZK5/WZ6Rbg0OIcWhnS63rNSWj
ZLUicd5old8ehDeRak6jGRyofOsiGoqNRvkvY4Gjokp22t/OxihOAMGea4gDMCERr3H6psXo6oFR
C6xqepjVw8AvsF/XhWfmefySLojHaP0u/qBuXWYCWO3MPjhKRYz5+AT1gZOaXjHzUJsXxxdaDMi1
6rzKZfHoYgcW6/8B4R78GnWjGFGMGiK0W03QEiEcmcJgwBNppVP/ndcYvFAgJ9v+EidoYRwco75+
FMcyPCQtcU/KGeXrxeZvORDJhiPKhtdIf+/49Lmt753oWprpj/SgN1eSFygv2yzu+imHqWg1ZXDY
LaEqXd59M/uo765uzkUrneAR+WcQJ+VVP6gcENJyk9AHIUhvo7J0SB4JpOVzPNee3AMiBpYOgvPp
iYXAqbXu1lIqGtoO+aMeXXOR+4bMioucVi+5a87geuuPuFQPs2EK6IyhoA+pvQhsq7/FI/f1RPK8
K8EgJCwFwqpKjB2STNVUztMxc8Z2hIfhd9LIMgeiNTpbocbR6XRQlEYu12ePTniwW+VaiMQMzDVx
U6mx4s7k7CEPwFFFBjidcFtTUEpb5jZ/34juVHmmHLEo9ZgfFjW7NwrxZOwq23yOi3IESKk0ZosQ
8H/Kyr8TygEyETodF+AyML3t1XFbhlCCawVv0nY5FFvb291uZCLEzTF5BAXulA7VH5ihsYWWfOJN
X3wPlLl5NUMCylKZcUy+2fNdyjTE69L5AT2iDT+CRXyWTzRQXsFzvaEkwszAGo6qEesALivrmMg3
fee/NU4PqMuEupyJoZvLeSPuWEJR9eoqBp2kUfnshhBHpJKD0xuI7CSCtT/YVsSWnL/f/74F16Qq
Fygxf9bKub5olmFYsvxKQdeOXYl3rKNY2jaB6nibCRMdtrOgdwMeMed+9Subt1TjNrWvb2lRzBFF
3mhjguBfWNUTn8jEM4RWZPfOme0Re7hFTfZNjs4vi0v0ZPysIlFeanyf2fPeYylrohDVajZeFwC7
vlE9WF2Yw6ID+3XB9vDuMgv4sBbJXxGQTpzV5FLO2TxuzzsD4ZTyd9vVFoE60j+ql63kzvt1qzuJ
U/6zaP0UG33RdfQCn5+vqLOEcJo6Q3NucrcxeZhJb/X45mQnskSgxKtFPi762gG8nKla36rFAnlg
J4LeRCxA0Ry2Txaz1TEGdp9+nEzqaxr9+Npm8x8sN+Ivtr9zStZinTWvedBH4JaCt5n2C91SJDah
2Sx8SwcNXZ4WrkZDBLaSIfmj1Xqoj9kHikyfalS5Y+gePeqoiabyz+6MkXVzA3EiwxbnxVrHAI97
tgbiko6pUeOu8PUNKtlzHJD+vwN5uwyqAgRbx+FCBRwI/bieX7sbKJ+yUmuhojH6ckHHvOKt++vt
BlfdCL6z0SG7TvZldmC/9n7v0o/WwzEFktUwICaojlHp4bRgNyQyMme8Uus4B3CZ3HNYzC/1ByX6
vegaFaFFAoBgnBaQk7OyhxK0lS5Xmkxf4lmgwEp7pgGCRELnOHFlU21HfLhsEkaCRCAMFnA89YKS
jZMYZy4OLKM5Aydii51A5UoocmZ96xiP5bt0jK2/i/fkCBayOWSCDDpHfhl0lQS78bd+h5iWhHaV
xd/b8etjmUkMGSKJqlMj21W6aj0sEKaZf9aWXptU6rg70eVmbZqV9o6k7sp5+mPO/krfovDJFBJs
NIw3E3S/dmQh4oCdvwILncW3vRgjwpZ5ed0j+fqrrWn+ic17z7eIR8xRVF361pn0oBFZtNzjeKg9
zq7DxibjfT6nCde7zqLIvlgEMcrxfFYY2pvh8TDOVlSUV+XUMZwcHNiVf/uzWY/ueZFzHLrdG19V
oz8trvJPnpGRoaMxJ2BR/HVY5HdbPYYxtzLADNOdPNUl1aQwprkuA4q1DVyOQLJTTbX8o5pYaVjn
joVzLBkRk0fiunBMbP9cyS4FwnpEIeNHM5dzzLsZhx17etW0x5uNzrNEDAHVNH6SWrmomsv9mm5r
XKPZpg2+Vl1SDgo5OhgSnutb/GtiLSjXqp9/EQpWeORCo1BlWZ9TYMSi597sxsZmHbT1C+mo1YmP
tPThby0fLAZhWRmV1r8z2bmQVR/5iZd+PBnwrrJo1coWpcFczJIJf/YbN1AzK7Nn0cNyo6FPQi9J
c716Hy4qOInsaJ17KUpJQ62IVreNyuP/3jicOy2XDeUEncTmkN5Yhb33CHtRoxBooAiH5HQDjwie
6bc/2RujspCP4ZQTXLCqD/s+N6tKv7JNEKjR4dKkL2IMTN65ljLT/X+TIgxi0J11MmLwZ7G4E1rS
EXUqj1xC1xS/p6/hi6d5mILayu2ZYgOIF8Svb1B779CgJq5a2Uody7RgHvVXIBrEMCdUeU8XG7rj
qOp3yULqWvXyaNFjEV5AQNDws+xREvfwXBcaJn591MRkm15Qbn/kI1h1m+tDMNWeonHzLUSsqJN3
kuGiyF4K1Tch0UZqCgthoNU6NXZjUaYjUqg2sVoDMINfrFbD0SjuOYyUO/OohVNKiYbOAhZZ0K1P
eL1/sNMA5DDBhpzBn+wSQpzCs9exLmqYdAlH0c88km96GtZO45LR3CbEKB5Y4fa66X7Sp1pQRrHH
97SEaeMLXsEEaCudSERcCq+RxglfyrxxSSxawL9kwDzFyJkowFmWHQG2j6AtxwZ5dMihzBVAsH1V
lT3oNVYsxo8sW3u25nh0YNLlVe/znMajiBqf36WRKUqtfpCkTQaxoN5SjFlfLxyMXMcNu4hBfX2Z
SCUQDx30jcGc8TLwOBY3h7jRa5uiGzm8S4oTAnCD6lp8PylKJNBH2s0WcQg9TCGtq5roor2LkxCS
kcpZPwsNKP85U/1Jn/B+N2HD+wzql8z8Su1HR4JEI6/P9M9fyCMRKsMkIWSsoAL+IeHKWYY1Mnw8
yfjYtFIVcPab4mdZfiFmsPWltAp8aLn1xo9rdrcUQprYWuIq4NyvbWU09R87KO0ofOj8IerFxNpR
BPA1OWyGeSCxjzhzwoCsYTPCq7zLxxGYEsNAGlOl27UfYHmhlaIO9KC8QGFwRMLx4HeL7THln/0u
T6DehyNuR9nnXEaVNMHs84PCh5oB2E2x7UCfpMSxo2VEaZq0kTxYq5YWtF4vG9H74Xk+vlS6QHBn
j/OUbBsBUjrqPpErNKvvpTnpCEUNMPKkeLD6m0h2AYwarEcJN/sRHvw2UkmKr5JAqaqxDO0eH/jq
LsurYC/+dOGx2n8hIyrtbfGcx/rynDFJE8afrGLgFNaknnWE/BroM4X7OM5mEcYZniFdvLg50rWh
zKE99e01lNSKGi6sV905MytJQA49A50Qd8s+m9YWHjj6KnyrQOP5lv2Q3o+D7vdXzyfvMZy6nwix
nnCr0uKvV/Amin9jIbr2d33AZIgmt6k+UCsCeWYikdewXpPoBboEaUoghxSYV4mrUwIycyS68GIC
8rMNqR/GIvMQcyAllR+FUPJNbx9BLVCerSa7KO3/5LJT4ZZ1uyYBqX5FxSonEoeOIDts+yIqzR04
mKfGAud9KUHmvJa3kmwW39XNr7b2T4KBBWvMFbcDK5yCectsbY8lUh9KF70lDlHnXYCMMW/LQKM8
vL+SL9kVWBZpY2Z5E+h15tZUhF0dWUn7afo8A225TJ+uxUGNx+3HJgD3DnjpglHdWOUW6USJM7kk
5cguqkWc3YDpU6M7+6PHKiAYVCTQy/gIWHdTdKD+PfMI58H+QGW/ipczCFw3BjUYHgZhg2u0Sgrl
fkrPUWSDt0pWwfR85bPts9RRwb0vsh+ScA0+bSDtUops+q08gxCJ3FqtM3ItZ/XxzXP0XBFuXX1H
YBIP18NV1xChGVjhw7U3o06P49Y6jyba872OFcOqvw4ubcbIm5dVukqQmtq7I3V+CAKLE9qt8gP4
k5E0rvX9Ssqk8Uwt9mwWGnWaLApyFlGz06S+cX2PzQKzdBeUI0CkMdO/ZPl2aOGKsJ4RpftEXa0/
b7SKOV0K0f1VTLp4vYcj1AHhKoY9INnCxGM39VuaYBZX20aaw0JRvZcJHEDKjATkoSUIIuw3fywq
hZ/+mFuE/zVH8khtEDp8jIgOy/d2YbXPcg0eWX9bq0NwlNHf6+47jEqZdZfcGtjGK3efrv/1ertV
+Irh6wUWsQVqgJXoCwz8pcf/0ExyGWeubkwQDLcvL7vJv+VNEz5SWFMny62t6zIaOREkuSXXFuD3
XzE5+yBVnrF1RscVdjZnxnKYakU6W4uR5lZ4//TzWa/zL7cNY7RFHvRJMjtiIoYIc2UNa0DmbIKR
mMrNi5k7/JBYpC4aIlfY7tNrcpPzN5dvk/SXxkD2pG9XKN+sM7n5XLi6kc2CIbLLl4UGoFJ5olMZ
uF4DPIUq4BnVgrwcMMW1oDzhVx1le9DGZiDGbnPBeR9Mw7GCWvRV05biz8y5XVmaMWO4BI4AsOPk
SxG1oFK8o5Dfs5MSBExtKEOmf/+Y4L8DPPtUACXk08InnK/NLzL02pMJbvDQkASIxTXW9Kv1ZhqS
Zz+fzeKZfyNJd9URHzRUWrPf4CtyVmGR16onp5Qxi7TAffBZWGCup8kfoCqbEQZmOX3iQjn/oCbd
yHkFftZ7XkDMiSCiG6+EVkf03X+kol06vPV9hrLSBz4xyQGiWBmPqO1UsARilLWHi3ymV10O3XDY
w9zDvBhy6qvj3UyDTphj6SZC7GL6sRnljqYaFCOCrBSc5xO7SYq8NREvYYFtqiORCgkY2kWVsO2k
AIAlTNsSetcoyF34ftqwwsvIzyvRKCyz61AKvttuVapKBQ6j9lQ9K+MdA1bSP2jhPXhW2ufX9+l8
hRBxvVTXaJH2yiD0/vzGpo5omiGK8aLEtghh7RFSp8WV+eZcL/CQvCyAKYcPRoin7B/OY+aU9G5A
e8bJ3nIzvWzVF8XFZOxUYT8UViN6k9yZ1mUHBnup7khkKj1O4T2VnU+tiS4H0kkadXuWojQAK4Nv
+jnipaH7BIF8FkAIRY0saArvESLH7D8PRirRUi/kSwKdKbzj+Z341YolSmAW0ExRJ7I6hTT2Wus9
UpogyxxQMaSSZeET7+MnM6hnZYbgglbDfVVrC7vX+4kR+4BQ1UpX61dxHHN/aHXwGbr21yJCoaQu
dkgKiKv6Xc+jnHf6cexg/THty9Gc0GuqsWx+5KwiSpZnT4wYcMrSIkLBLgKQUaRQfS4UCr/SKow8
PWEQnpx5igNh1f/iGgv4Jl83mRbK7z4bF0PTtBmnno1fv/HCsk/TTt3r+2PX0nQl8QR4lcrJ7hNA
HtKLVV+I5h7jWQxjBI34YmT4Yaz2gOLMg6yh5/KUg8uPuUfeVWOUyGx9A1320KyQiK/nlzb4hO6Z
4JuYIC2DxhpCsks8GLqfeXOkvyafjtE9/5/yWwxFuDjOzgutN7mefptANbzb+scfRLCpDlFBCibi
O++EIpGrIsqLNqmyEILvz5rhjx9t12jx5yc7YPUKZ4FUoWm88Z/13r/d315ZxS6TtYZX5a3uz6Dx
iCt+5pskpCNbhrgdutAW/kjBwWQpxmHSrsUAbW8i620zA68RW0lHN9WBG4yxaz7MfnQldTjUyx5w
zLozrHMc6ZU3XCIj0VNW40XCwqHEzuOZOQ2mSyStKsz808cXcnsRg65mMBQHzHY0X5sukk5RTFDM
QDD2La0hBdTvKnyDSSbeqnvtrN/orlHejx9of05333zeYz1Y6vs5AZLXBYV+Bee2ElebUPJYqyEf
QzvLGufswq57Zea+Ku686jVGROWwdOEvmMI0CqK5+HP7NcE1mNZXlYAMRAfG1NiM4ZPiyw9OZ6ns
EDhQTPcX/aKExK/T+8Dh8DZoLx4Bc6xBFRhnj2Ju95hG+41uomxI2xzMRdGF4JI0mr64sZm+2koS
zFZvohye41MnDflfgyex7dMVyXyffMpPTPH+h5uonTUxY/YSBDxQLwQslA+clj+7yCR8vU6/qU8N
eX6rBUdEgYm0qapSFLS4Zo9oIhEAYq+3cZMVVoI9QmC9S8JnjpzVVNiZtqQtBZZsMzn7ri/sCtS6
F9whJQElu2J2FiGDLaEzy/QpzKkThUa4Wz2lYI+EGPGJhD0Wjx4IyyXyP/fR3gPIYzWFEM/nEtIa
FKYLlAtN0y2pMxps0N2bWTOphkN1Nn8fDa3pbUCb64mMlK+6lNcly8GmcR68uRWejtlAQ1huaIRC
TowpK9fDjEUJCmd3wpbWEMK9I8MWliAZdsBtI1xGk0bcYNF5IbSo/KOHVzsIW3oNPiwP1Hm5ePzo
AU+G/37nTdQuHSRAx8LWEtbJ5nqPTQLvY/Y2Eco+mRVsyrwLrNh3XNkNACZKiswg08vrpakPqmqc
vwvDV/FuLI27tRTtB7NGYYUjhYxUp3KhH789aaG8xrkE6hqh1yYm5243f/QdWfAQP/HXbYJwYnhe
dQ3amZtJSxFUqjOx4T1U6+uGfaW0HZXiIp+oieavB6lpPMGE45BL3pxS9wL4G3kax2vIdmGc+U6j
CFqSWywDb450cxUdKhiFzs/SLMmvJbewcPOSQaAXo4VvvR7CyMQKbODXRXJetGUCJ87ZVBwaFlCa
uh6VxC/pP00emT0szIJJaf3YgYTJRF18dA88dR5ZfCPDw2rM6ZVOhjnMzqfX1eHf5Nk1V47cGlCp
bPBTDnr6qzabdGlJ1ZIH6asahEB/trlX/9gQ9Pp4aO6AMXP0xkmtHV45VDGy8MVzbpWFhYv2611X
r9+rJqLJ2fKN9cAf064RWG4U5mhJ8B+MD2e7AxXChsrLGk8z4pbNU+54bmO9SBDH6F8YEAZ6XJ28
TUmP+3sNv+GuUj6YA4GK7w/8cfQR6l+uP1eosarjoyUJ9R8gXeajg4xEG7YHDtEocLOX2CZEsGb6
FficGvel/sdfKOyhnzpU9H68A/RZFGTL1awiujNyULsE6e2gPY7QANp9CZX7TO3a8dNkh/onoa8o
IjcOv1lzac3fpctmZX6OSh9Pv11iJbNdvjpuBYpV735v+KI91AAHd54Neu68U5M1al9LZNUyz+Kn
TZyJkNN+7MLZxLJrifq8b8ifhlDuKSfgoFtlIyb47P861ECbR2xqlEYTbt+6xQnXaA56qtgYeNj6
lYjn42osi1fT9iJ1MOOYasWSLiUNAziL1FjoZ7CJqB9j5GqP+OOW0rXNHRxjxpRjXgYxWzoDqyAa
/J2Qt4tWqncFimuvtrngfRTxSoNZYe0U5vSxwFnwHftobYEnT4SfB4gQ23G/Ke0lEoF42hcWccqp
kFO5HocspE2iExsashGyC7tHGUy0F/C2JlYUPdtLzXqYTRa5pSint+xIihAYQMGEixgbyySCd/28
wrV4jZTNKBqW01BQg5rhTpr7rOl3AB4cJqzn3vHNWsC0O4A7lze6Kv7meMu+4l+EBxTU6BlfFGih
/TiiiqLTikzylwlI4O+oCvvTS+Vf6QXGawLxZUe8Tn9zZvkNt5rB5wzy08z0Y14VfVJ6FXJuCJmO
rDXizA8LLr8QfEmztQcIl0gaqZCGwvdxgIhsDO/pRPrgsr29wpN33vjWjIyVsxJ71rmFZ4yw1yAI
S50WbPMLTCXerbFCPjMdf0NlnBymL21REHKFklfxx7fOfWC2RWBMtQaDb/F9MlraYcD2C+itojjs
nqrqAdRNPeMCuwnmY/+hEz6blAv41XOteEqUhp5dJjoYCuTkaGZlSiq/vr7hd4sdKPTwVYsZ+wv6
AF/UNbfaw1YQ3eBV393H4NoycSS6dFHQy0/UXnSlCD12rRDRSDskosYBRdRRT73wTAh2X11r3kbe
+P4bg73txndfGqaERAZga72Quh7uLU1I3cBkPqa+lZVGcH17+0Esd9O4QTOMhp4YsZq7G0eH4R6B
KXcAjsADUx1xXgYq81l+6d+LK4Y9b8WWMxlw6+CjLh14ZtIUtI7bi8QCCPiHcYknXMCZMVMUGscO
pMD6BL0KwF4bfNYumb6t9ShKkjBXw77g5JKhva9m7yCCfLdbzHXF++jbH0tHXFpqpkYiIfCUpkRm
w0ifBPQnM8X0gdyLQxkcYl2zoogWSavroUZkU/NNt5LTO93r645Tl9D3n05ZKegHSCSDDZTkdYEh
eUMa47zh1NbvhmAZL1xOOey95bRpKfjacgnZXHHH8YNxmbaO/jywGU9lygccgow7R/YV3O8QpAj5
KLXzgPlDQPucVq749xbVUPPVQbQX0tndEza53xLGUvuZmoxXgVJ6Yw4df4DRQJkYAzzvYlT48v6x
WumzA9VHFD7CSMU+v6fY5txTTw043O9DulYdkaOi+kyV0U4Azg/M7PsAIfsLhL4hocbW+Gk1ndGm
f4d5s92Dp4/ghQCTRY68WShQt7zEeJsrf9dOw9zz/tB38UV7xKue3PDHn8f2FrqE08i1hIOfBouO
cQgEjHupZjm5jI65VNeyMK8PzzCyiKp2bXSBqtPzMOYNQ8EqEQ5QVEhi3ukk040gE7KKlg2jXjdW
1dAC77LNv4HG5GKi6PXptnPR73B+4bM8LjGkfejlMggI8JB6FKllfCqEZv5V8FZUUtY4xWHp9wSZ
TldX1/XLZjhoW7fZiTUmlQtImwWSuz39qTLonMXHFtf8vT88Pq9XcvLzWTh1vow2idsYyzIFqDtN
BBlYy7T/DMNX381n04u2qaeD7VvQcjyPSeQAOON6c5avkKtcwKOGKMxLxknbntCaH6PMBbZPof8e
tFdLz2EXJV9yiQ2MHVnPvmM6ej9aG8YP3LLD+Z1+cK3vUUfQSivMw/Rp0KYIuNz/ppM4r+yYJ0KD
fBI/Jfp+XDCJ/1yyUf60XAfLy7WJaDgJ4W2tlbs9WmI7/DLkwxzD0dxwvtrzY6B64ztceIRQzM5v
ATyJA81j5uxDbspdVDaM/LdVU9yStBwaR6McYnipSOWCiZUjomzkNZL9izOkCt5mQpYrvjK4QJBx
4oCdZW9mP3v7b5Fei61oMgOOr2AZAM1uBFzQAW7bcx0V/gO9cm4IxJXGVfSv+GY/0UD3yWqIkl4F
jQW0stvsy7Rq/UnFFXJFJWHHYVWQOPTp5Z2D2SVVSMiXPgoKaOflzO98es261d3gW/vMfoz1uGg0
apZ0WIuhYc2DtQEe+q+ULgF5L1lGkBqwoDLCsQCGon0livHg8nY4PE5a6WYvPSxzAx4R0CURNJ3A
yLJ6dh0xTHuT0cWGpZm57TF3xf4nti06ICed0X9KZi4rhICUXkPWcxpJicxB2QRnvHZohAaKfiDA
p5/enFiIdjjpSu5WO2BRyU1tSaiGv94IoyhgPiQeUgt1o2eSm5vYa0On59zVIUwUbwNvie1aZ+EM
m3B1jw7S4aRuzXzTN8q9m+ji++vBs5JlMb7rsnUduF+u8FtXxBbj51/RbLZoRZSeoSYDpa20P6/5
Gf5mpW1bPtB2Qg5p+mCUYQC5g0QDkVgtv8eGUu05Zwg9GaT3uKm1JjaZ2CfbhaCRRe/MQFqw2JzI
YUGJz+oh5hz4S0lssGKWhT1B+8Yy3S9txR4zemIH0Mmln0SspjYwmHpcYuwilltsrMD32FCR2EFQ
tVABgTF7H12Cavxz6FyTgMojyUhO0YolPjUyh8GpFLqtzlIT74b8mOvnOyTaMdVtBgwnc+pNdUPU
ye7h1LVcC5G13PTolYEmvOk0YVoPEJgY2MEu3BqnQHnmBm3CK7p6t+mK18SGyVn45IcQWuAgyTTL
W5TryYqIQSsDt2MyBRj6SsGbwp7kzHYfM6RxdxmTlPXiOmuM++5bFCoZ/KAdt7O/msOqgcmfy6+G
hGSHi8ByVS1RjyY9vmg4zYDwGohtjqUz6SaAAG5+RNQFnEfjn0yc4KJ3aq++t6g7Xoxx/n1hypR0
twCEbD+9rg1v1gamxjkNvJ+d70O9EExiGcCwDjvoj84MEucfLvCgWgRZHIbTj988iXErPDOr1lC0
RwYx/TLh5aJxB8ATdEEKXhCwlIfjCck9Mil+iAdFvvNvV8t++oupKIi5UPbvhT0VC2VnIviNEWhG
w9HkLHlyoxP+a9Yl2Erd1340Ih+5hdPjiTpQaSxIl7E8FGgGXbxYDOJ44ZNX50eI4fswtWdaaoaA
EmyFBqzwV0QxcLDrucNeL800Lv6diXUv7GBXz/pmtSdC1ffOUU7/MdFfjgYJBCmuvFxVvznywXGl
Taddfm5TUnvPYhcPhJ0hnWrssAaJzqqvIXNXmyRF4ILpGRYS+m9xctshM0bLSaME62ZBwmxIe8FX
KDXD+YjUjwUkuHeWzs3SWJ5GpZ5jWueXl9mAMulg8hLNXuNaLlWzIaLrzwErYAJvXWmKCi/yuby1
dJVZP1LJSqEj8N4Uv+aiDsY7Hjfdj3UdDHhC1XYN7sZZLHGPhNMsnOhDd7jbBskvzTKPySt/I9wH
A8+ktKEAQtWfJ+RdGmG3Thl7YcPu7U9KrK+NTuAThsuBVf7e/ZF87feKxd0EmeUsnLKQQCfwQx0e
cw44wxGCpaf+bgc6cuaX3FmCzOq5gJo+RD8KpA5vvPVq5IHyY4KII3g9ICC68PW67yvFjSfX1eGZ
wqPCDx452kAEgu0mUE8Ulx9n8Rqyx1xRvPnB3WfP+mcKXm7xApu8h5QPH4W3oyHlFyPjRiNn8cEH
H59Cr2mDYyWR68xNaxvUR1tb4jlJcrSINymhnKcGVxjfBzTXkyjZ4AfD7+u5BfxsHCtkZ+hr7iJZ
AFgadBEWi+6f42SSsmYd2tX6Kl8m/VJzNsPFYkrGdsbZh8TMjqtRfCQmonnws+4t9r+ZaJF2fFOz
r3csV7p5m/xEy7OT8WsCUCP3eHjA11kuUpvCK/qeFGDebg13HxgKKRYSfEjufN0EjnusjCe4lALj
iAuXJekQz231SQOE/2SnV1w18c7m1Esw5TcfsqZPbgqmDBKan9nCEtlm8CadT/yLwTEbdXkSdCj/
5I8gqLnXbqbfQxDd7cZqtRHRi+G/gGCvK5j6EGWuqPPNcoVjhZKLhgrj6QRtDUtnh0dF39MLEjzF
JEQ8VvEl7zuqIDHa6ph+LWABqsg+OA3qhR+GrinR1XtvowDEwFd0nupWwXnHtcISSfNyg6T0CpGB
8NZWsXIL8lBharFGGJTSDCASk7lUleodxVE4s6PBrd0QclYYCwEsB2Fx1xrfn9bZs8J6/m0/ZpyQ
pKADV18PLH/V+J2eKzjgde8RzQOuZN7uuGHMTS9MUaT3jPvcauBcTjNM+jeOQsF/VNT54i8Ke7r6
EXjWpyP/CJuG0FS5WQgRdV33vxZchS7ec6mfEpg8viAENK1ay2j1ASgAce0PIKoz6j0yPcoCjcT5
k8PC6iA7srD6pfBYxSuuodthFP/I0Fb8bwV/qJhF63BJ2ucRWbRYkWlWjCGiHy9XKz9I3uIvCHqI
6EDKdgvfrNqsFCVV8RlQ7y6fxeUdmYbi4/vGlYgcxX5vFepwMHEXzhaFLj09Vr8FJfKrNiLzMuHC
poKo7eAgV1CS2ipcEZ+PAMGOXm6VayfXQZLZ/djVAoxQJw7c1yx2vTOnugVaHPQE4eTiHOnSmBPX
owLEwgkrvoQ3FxN8/13KAdBMekAoGj5FKK+m7OKbdhDFwjOaUCIe4UQfNvc35Q5BoPXsq3cMiDbX
XeGpotVeZwp3zbVTpBPi5V4jTtFuyCUCp3LFVjelEzksW+I1/5Iqug6QP6UPMqByGv9DXFlBtWs+
YtRov2WXArVnfuNNEzA21QGVXUc/M3ISVA4P+bElEEzOMIy9M4kEDKpMydPlwRdkr/OojTLB8MiJ
uWBIaSLMQfC3OM86kUBubMz1NKA2CCWp5oV9bu3cIjNH3mw/1b8B27TnM12iJOWiSv7X4ejdkA5j
aiGEr8o5k45vPpWRN5MIOroG8EA0GD7pVwQFWxf66o/J4EfbePZFprwHDms8MRkWCXyraj5AQYDz
hy50eSTF7HVuPBfHRsQ+FmQ3hkrU7y6hb4zlbjX+tA04V6Hdmp9Bq994mUAygHoW264+EgrvG1Hp
VRj2UUVvrXZjnM0u4qKhFiedfbjc+Hmxna/CbUMGGbN+cpQErPVW4QWNRZmxAXXFUpmkpEF4thld
/UquXLrGycOBikXDMvXgOQ4iJNpWCVPES5aWda5xtrAAJsPIk7Rmr9U3mxgBtWP4tzqAZcqdniP9
z5NETZdIo64iv0e7AH6WfuMjdIUf/ZV9NmNjh8BNUv/PnhxippT/fjBYkktw6+MhzOyEcK/1TEk1
qa0tjzxVFqf+nTMe5X+mRrOG3+wNtJqWtg1bTdGbllNpcB3YduKLTE8v1KPxJq/pQiB5aObE8Azi
JQEg+Eeq254qaSSkUaKYVMhfoKIoor5FLWe07/EHuk1bemjX7jOckjS1wcuG8GkpwxDtdoseq8x6
1K3Q69MlFPAZ++NU+zXQEmHO5gFvckp0QLIU8u18VLiH3/zQmb81AMtHyjRqHhGTKdu3+tCBC3A+
TSKmyDb7VxnzjroLGyGLLO4LSpCDyR7R8Cy6mLKDT7NZ2e9jrPWVyWfqUOI5pqOleisyfOcPgZXJ
HZaEbyVx7VDgPd9Pq19UZBVyp8BAuEsLmnqYDxw/kizTbPmHFXZcOVGqNm3pNH2FxDNxtWAA3yig
sLnuAMS/Yw/Su7D3CTxoQZUaB6BRHwjFKJk1HhC9COgbPJ694cFYNSDF4Xsv0pp2ne93FDP0zgf9
Ywq1nq0EL4HNLgQffSwd4UlYNSNPsJz85OpQ5+S8mVhVksCzj/Cjfxk5H5+WEgNTST+Cu7xqzU/B
uRwqn9wywBTenx++7+pAup1fcBlNmE7n4f2dX1eN+JQg6/tW4HbNs03u+NNYCmJYH4Xhty3oxTYw
fEhDee0SiXBfKKl5IC7onr4USYNcudNIc6WXoD+fxqSi7DvuFNrcV5kC+WW6e6s91CcxGnNrL6OL
9y0tfy70oc3JY/Aw2j3O9cYeViQdqmXk6RzLikiW2QhnZh2E+aqMb0EOuJFRQTOCdUEATpuQEF/+
mw3w5vbijU5n2BpffkeITn+SVe00r8aoo6BjhzHGeoyh5giUdKwbDssNDHhptLboUsr+8UDb+RRQ
zFTmBW7XWaWFGzRDfny47xKssupBrJLO4bGzTd3+k4K06Hvc5hLl5WcQIAQfV2BAaqpglilwHvWa
jXICXAu7MR9flVDi8hyq4qKWGLJvBDQQkopKOwke548niAQAhDi1kTnCPgoMT+Zlr1UJaZysbJPV
n+v26iixb07zeoRAucHrkLaQFyi/ntJHzJq9jCdwiwjDx2JVt0S3E7FjsMx1uSsq/tsJzac/UUP3
qKL3HRfTq71UXl6r4dfsqH1QhqRWmidPWrLrw2JdruM9Ehi3KPV8I+tKeon63k1DvOov6smELc4d
ypBUe2CZXsYuTDqcGx0fTKPKvaXGtSwXTcGW2nu3QfaPEhO57nMRkKiYxT3IWJ95Ry8Obbxn0n99
UrbZ4Xg8cSUUhOEK4IVITNvMAlsLxhXuk/cYIArdlcgOwfIaeHZ6yWJt0b/+rmQvJKOqUe8Iky1I
OHeV5UDq+n6dF9DRQrjXOecQ5tc7nLTtOAiS9Thsrbow0BahKcaH5UhgBcIUR0j0t2OmS5w71SV5
gDHAseeUXW7XlBsNfOfdra7/iVAI4iz4kwtICAs4n8xx14nI1lSKUJYflA/9Omp8cjFXIzd71fRw
iRWsxkzcyvyvIRNqMLb/q8rGVleam6o9EJKwGqSYeHp3odxGPWBbyraCLo5zLmBWo6hl/wuVhoLg
qNK6FtEakzyUCBrTrNgZMMAsvaoJX1W/ylrDmGTvVO3LmhaiTGtOp12zO4mdJUAVtBVyrs18JIPx
3kCnMY/rOnSHQMYtoSN6xfI6wBwn15QPhlmO5/EsIY2u0kiVl7CpF+QDX0AcrkZ/3WT3AHZAt5PD
k0L98j5K1XPqGDOnmo/agR9PuoFecM7sp2ejvwBI+GMAl8DsCCalUge9dPrsg7iY9oYw9Z9lvIJa
QqWwXmmzq+MUGhshDTLwpu6GJKahuMm+/pHxZIsrkKFFzqbivGrpxXx974sik9Mby+GoHL/QXsa3
UZnfuu00XvgxXIR7zzHdELHCLqQ3q9c32/1mvwOpwLUsVi8xa8kiQ10j5M54oFS1Aca0mLy8I1BU
b/wia+v/nKe//VMXKXUCWkv5JlC0vRgI+kYLE17FVF63cxOPDR2iHFCwvgwPyCnNcna7Kwbhevaw
hINFjnIho8Ikk7O+Br4xvwN7jHFcrYD6c+qYT3RK9B5KXJckp66dESIB3ikPrZg48S5wUp8X5yx0
0y9kU35U+e810c6Kwmil4hn3/FaBHz6XQK+4XVy6IaAHNcWuwOjQSXhfk9ur+Crx+bt97cyb5Le+
YpLQ/ovxVZ+8Uz9iFMqUbg1Kt9+RRNYrs8v0Y+Qcwyg6eZHz5ptgYmQdBgecv6tBFH1cUofwC+0H
XuC66ePYwg+lOOidwqJEJzIzTVjAtas0yWRvvipAdKZjq80otVGiQTg02UY3dwsEm/+y8HKjMyMH
q5KBesJVjPZOnfPqd1cxwmB6iIBhxQDmWb6rU3Uf5PEh6OxXcAzR5PjZXe5Qv0XQYf1L7Qp873ia
cKTikh+3iUtZNPmuCiTXV1wQtv+ybmGIQ1Aa6N928eNZiCSUBgM4KwAmNYdsYg9GRbSZfuTGW5OI
BD+H2i4y4IrUDJoCL1DMHE9Rv0/qVhfTBC1/2BcY+vr0vG93esNfSnrvDGj0GJx6y2BU9WwsjSp0
o25Hh6wDA1avszxBu0PB1nS1ZP24PJl/6SunIzH0HFNidQ4OFsr51guZSEBDUzvjRDzIOlVOHoIo
zchCWfVET4E8y5+7TWJS4IKyp/nloBk3j7Lf7DQ9Rvsg5EXwa38hv2hXJUgGjm4yJeVM2CLiLQoY
3n83QwsmGp3qm+0LgjT2m6cBRP+716XqY0+lGEJ/Li0an5UIRQtoM8nLV3+m7K40hEehOX0l9/kI
+zgnS7f+WaT0AQ0LlpPwe8gSPJPCiP444l/oyMmllWBYYiPStCIiosRb0MOWEBiaGSPGeYUvcQJT
cmk/wk05ZpW3V7zEt/a5NlnepRKbqUDOnvLK9z+oTR2et9r3Z8jwzg4HJyC1VnG2p+xsAhyX2rL+
0N+fC+YgnRyfvq9nIJbK8ZP1wBR2BIc2CBtqWDUQH9ckj6JxJP1/X4SDtIo5OcBqFMS9Gk/n/mEv
e3NM7ERqVGSCIIJaMBjgo8mr/VMIlERqC/zc936Si192UJi0yJ3oNN6aGHN9vwM9m1k4OSQVpgju
+5tGbVnOFhkjj1WM4SDcL7raBGnGIzND2wOQ8Sc3eIa5fnTsTeImCN6Hil1uycGhaYsITW09kAMD
OvPXMcMDjXqXAPnD7BwLgYc2/qwRcQGkNPIrwJpuV8IakWqtsYwGwFv2K8pyiIFdKVHc7LzuHo/J
g7dBzpi3eabiE1gZI8LmFolXOwy6r20XFyb8y0s/17ykRST9cVt5WoFdg4MubBHiXuYNvI1+9ELy
5NRAeTsfPgposxXQ36lUd0E7REMUVbAceSf0InVSRI20oHY+ZF4zKu4Ns0YNSzFffRIsOv2lS8EX
shfNbTNZ7LWxIPpT16wNdAlf4syPF+vcTHDIdJGCsdUCiQk/2JcFUKPmt/VP/nbGu35DHNg8+QX6
ruEDrJIFvUcrS+BAU3bgenjh5F88+xI7RMHeDkD/yzPGZ8047JVIOjpyqwDwOUN+jqxN46D7G+sr
t4YzEHXK5h/LfRobR9AJNFU7v8i/50lfNefb5ohP8viMLjfDohQBlfxnGSSiZXvNY7SxGtg7GmdH
PaPSyLLamEaArk403uyzrj4FH055C7wQaYxPELzX55BqlIa3rvNQiVVRg5oOiKTJZIP7HO2ezdyC
dVVbU7HzYZ5s9ePVk3k0/LDQYkMEkc6N2z7bNL5Of6oqD0dZrSHWHuiwFQfWwrHBLhlhowT8vVxL
M9m3n3DkLnwoKnVR9C/CuTjjunSklIYzlp0hhyq4+v7wXIGl+TM+wEqorGQtS4e3Vi7ytSdohFt5
auI4Q4J7cq+9gXqGPA7w+n+XN1O7TXsiO3XBEwxREf4aB/NsI0MntAVhYQARQcI425+7ZOKtBcOK
PIg1XH4LkFYnUke4razPTIjvA8Uolw3kFPhCCpm1lK8i1gmuubmG4pRff13ZjzQUxzhoSPhcAi5+
FgJuN+YMH1CwYopi4Wjt3TMSSKBkOV02AROAr6/rLCTyHOxMoLngGtDUhfsjMKgWi2ikuIT1ZQMq
Y/i59HnU1z8GvWqhwVT0Ln3OO7PY+xMNsPyKEHsnS40dxms69uvuSw1ZNzNLLgmjPGULq/msLgTy
DypeNZbxpKj9A15vZKY+UNu+dhgpoDHww+xT/Y2B/cRiZdvDBeWf3g/uixdm0xVAO7jFYfcb1w07
2VOJy0G8C9I9Tbijr9Kh3a1sF8dKnxTktLLEB0qGIDLihSGeXn2PiR3sla2FTyE1vZXdka2IQjwP
xF5TztxyuIm6ZjkBSe0jOyxhvB3FgKur1jsMBOldtuby5HHx/i9Bi2C6v609x2jYqqvHhR16VrZG
kTK2b9MpJIyM6mg49vK0E7BeT8nuDn8D+t74q87g9mEAbqvMikZjRshqCTrmGb6fwA1+NJdsacI9
kxf6Eu6hanimiBA17LqKdMOEBQdZ3IQIGaAzBOpJNh2tILLDqBICbsO19T6JXyQ8iXMY/rVi+yya
q4zDvHzNx2l8x8gZS2elOljv3kmZgnCcToL8VpiRkHYnEWc+6EFUNnbI0Lse/o+kohNc+ykE3RVA
3Z9h2EnmdAHqaj2NncbLH/G6T1feh+czH1nmlEmmkjwkga58eBMJyw5TZ084RgFGWzpt+2132qDL
tR8D/zkf1GNUV19n+JiNo56xfJ0yvL3Vno06gM9xod1ajKqYCllX+J+YDs0H/HddLmtyGPki5+OQ
M7XLHptoTKf9qFNHWa3Ad7HzK+ISH8RinqUqs0TAbbZls9PaIwfeGVNhnTFmbd6tXQGziOIYKMh8
TEJoGg/j7+wHfmLb/PRtDCfZyFc/w0VOZbV5ycR+kQfg8eJJ8aD9Ow/pAwA5zONSJk2u7fI3NiBx
Hb57nln2OaG0Wz4q6wnGhaTZp2DyjSQrGEZDoej2obvKIEpk4vEFN6QCzNhdLbm5UqSwxkfM5c7k
Na4pbiRAd8HArcetzSF9zKd+czyZyl7V2/UIup60Tiqk/m+DbpuSW9yjWS3ofhQLoBQ85qVvdHeR
hEA4n4+LkT4mHsJcjbsAoC5aXF25DrlauUYFKqBWgJQHjDoCDWeaIMTr8OlwzEb4/hxg92pXVyYY
gPTVz0ZdhD3ConiXlaBB4MgXenEqwV7c6K3OIu62JZU8pGLQzKNRNknj8TRL+bpmtl9xvZdZDi78
N/wqrGVQa7Hy1mX7yZyIH4AVWI7cF1tfluGcjYC5UD7Txw/j08IC66hIcZAwLr5IOzF6YbTtuqp7
SoByN+as4dqr1DOKAOPAUBtlwKJ2b71EcbC/PyZta3HEZShHrEj3PQlIEYSasZSc8S5baPxTvTmV
APAAMTiopT0cJ28MKDRV+P/gpddlpImwFh39Q5LDym9/Ab3p/2VnvnDuoU900KbbOmuMwzJ1nVOd
raE59G99lVcaG1wtx9MY9UB5VanP/UBdjexfWG+wcCRDdVSXmzvwyEIw3sGL1mrWqO148H7KpPXV
wcoJ/khqR911NeRbeUHLggXoUQF+C+wdcoTn4tHykQX0LsR7AmQ8kiJV1je2PYbmzqsFVYW0PzPy
85UCo203BtaVB2YdVXBDBM4S+hrANgyGlFyekdgZuORRqq0BFrZZxLEU211C7kMEt3goa1GVUSzM
XMKd+ei2oKDcKp5FSzPERGtm/0kwAe2jVWrRmXM37EHgsONkVoXdHGbIbPOgqrtILUaMowlDZa3F
en28ceJYF4lOxU1HEm8kSWfLP+AYSt7kxQknLNGPkSEZ05TmP/uDh6gM8aCqNTHoaBSjWEEvw/fz
Nd3Wl5J9CdnrVZHDXKCOVUD3UCKtom/Pu0/WKWh0pM63X+y57kSzw0YEPHBITam9364o61E/DS32
w8djPJnx4Al4bGnuShE6Y9QH9Z97G9vj6ITzMSnasQXPDy7FNRzk0MAcUZy7gvnEJXUddY1x5yRE
3nJdlyktmnBaXY9kv+vG49YgAGByWs7mk6VPueZXWz6kENaTkItSOSYi6LMCbkQhQdv0hhl5MoFM
A9mBLxBKNN+Yj5L5tU/5mR5uUVTGJYBkgL9BnAaK2w3E+4i5GEG7nzwsNs5I96h1pmLR6eMDYmdL
2DBspBhs6jzX6j0D+rx4rLbF11hKHS/rGVKpQGBAwfiYGJDRtYl8dnrNh2K3QL681Ui842lS2zbv
BcMAR/5y66Y/30p9lZYwIN5YXEXEcVM8J4mQI/kEe8OQXkVj+qbquMMwqChkEXrBthwG10fopWJA
vNEsvlKLlLlzApkfZd8b2A3tyIpyOK+MiD2LR/gmk8akgywl7v0tjd/MApRg6TbXie3lQeG5AgzG
7iveqOMBWYQlrp1aAj7i1Qoaeo7oOmtfd+wMMwkLVuVa+Ce9i4ejry+WVKqtdLxmyzvx2Jz8xfU6
KTca6bHHWKkcwvzcX8B1ePd4BteiozDYzhr0/cWpMw0UEFT3dolaQ5kLe44DpZwt1JOpqoI4Hk2Z
3vlLQGIII36XI1+eD2HvBAVjCkI0TYJgRAdtR/gGYM5tdXRnATvgaTuPzhWFgrqWvdKolNXEb9QE
XQSxLk6DwuwB6WCpVmZhqEtinV7Obnb3HdFeLKMprXkk8FfwrLpPkILJJp7Wf+0M4upJajfGL05q
15QZ45HYlPXhbz0Dt9w6ptE70mmrZCI9h6uv5xoyQaCWIyc8F1r2D0zmIhM9eFHVhr2VVa0/md8X
LiXGuaByRtCqG/pOSi45fows7+C0UWOutHFjakJgFLEVhsa4feEjBumqtI44B+kNHhOp+RieMxc2
iHJ3g8b8fnwlYHhnOFyK8vNe5QAyEGv+K9SjUD/jCMhq+77dNlQswrQn9Cub5HL/MInit7P3EUew
Cv3iRHvVIINN7AXe5IRAe6s1Sdj2WT9xW9L8hRcYcg7OVPBc42HG2sXmSVy2Xpy9rCtaav8y5BXH
+8RBuYli/POfSO2CyNKHlkTcb5RhtT06Hg7+NXPAnUJIr3tDSTuzzLzKaKhiMG+LR9+SuQB8KDqu
gY9gmvotcrfHMdFlq3ynmhChtmQ70k9ZkCEcp7iYv6Jr0hTDFGtLW8g06hvlSaSyxBbjx7mj8B3U
cGNhnxpxawShnzeerKZFYbE+J2/Uf/CdTYpaX9w+Phj/dvmW8IIM2JKJ4m3C0g83e9YQqlES1g/N
fQveyNhW227ZrXdWKe+GQpR5BAYz9CqDU2cMdqT5RY/f70BnCklkh1jrqepuxK/3F16PZ8RUtEpU
lykrq8us20wP1PaIb2cj9ePon30QWLQsFnUuJoxy1pVIOvZQeY3RTwtqLbAd+zcF4OTHBbZv74Gg
JrGSqBut+ZHK7Zym7QhgtVDeOwfl4lD+NC/g4vFqvoWf7lJjyV8p/Fd9SPPabrGrTUE8N+AtW27o
RUwDijf1cEW2+KdjCjymGool0fU0ISQb7Qt4CJF8wPBgMNq/xW4IcZHlhR79KweYOajinme3rY+n
RnAUlcWSr3Xwqo0zC5mJTjJrXEhuph51yV0aIzVCJalUt6sBMPafWazR9O/r7HskVB5GdKFEwHVV
6ZAumGYvtUH6364SeboFY9yaYAsgjqxua41l82rkTiObsUsR4Tkeah6g8hlJNq/COhObde3kJ4Ih
pF6jfuJL/H2OCsX39c6KZHxOsPsljdyweKYkvWLeT8q1fIazvtjes+BUZjWt6yrYHuXJyewf/sE+
oTgY0ZznyOejVPzeK2DcnGbrZy1B9fYAT7zWBsghB9ERVbnSzZhHHw5UrZGGzJ/NJK34Za7UnhjX
MtAKhpurR4CgDiGuss/j2pQPNNd7Tw+31bm84CabJu/FsDc+4GB50Kw1WtS7SpjEox04d1ugGdQk
JcX09qgDlL6vqc0/Zgw31YEDkPFNpQge2xwOpo2QcCUYMrzSZ7bAdcM1RL64G3S3Gd6n1oR4ZyBm
5HU5uvAlwHTxZCUlMg8vTfUGXOCJh6Tf+uNRVTYXv81WUXT6cMJsnIn2jlpGYzCU1JQasGEUs/gb
2237+4ycIfgMlZx5fuUMRrGNYx2xihdN7MJKhUk9Ysuhiz8/TbXPNwDD7/IGILL/YDceqjDoRxFH
6gSQoD9rMkT9RvLO0DlfndrOzd7oOGfUVcQRvVpO2IyU0gnJBfHjPpQt2/goKF3m7ZlKykESg7iu
rJuYK1nM6PfMLzLoNAdz4PESr4njC8Ekx3DuGD4b6kXdEoXcWy4tgPyJxIH9hHI3tXh+Ul4DGQGX
2Z9HzBdEoNVWZi3KZ3jzMewsjB2Ilsjhu2aZ7oL0S7vNipTvCMTGqsZ+9jPJlBuaqEyZyZ+lVdrZ
BXbbc7ZUrMmhIlleSQIJR0Xjy2Ywi8nLLxv6STuaF39i/o/t0P0hneC42KEj307b03oHvXFzkIyo
uARxl4PbCwtZj/m0FMYwMIEyInH6FmXtJ/lE3XOh3Rpyc17zKGgfyZ4IH55QJEcLxM+oebKDeyg+
DJ30kkcaxeuFq45Ei/qmHkWJmwu5geIKCacNS7PNl/VRtuPR1GZl/LCtCPu2Bn9Auv3XOwaopyJS
Af5V+FjdNVwEZJR5sigAH9FjmkJxkunVo2i7SfEY3h8q0jWAMMRCoQTea4UzNJYIQk0dGIP/8aLg
HBis8oZgtDFJHfAh3VdWPGHWI1dtP9DX8PwZ/CayXIfkFLasXn3lr/4HVElryaLI5DBoLkYXXXqO
vNfLw0BJc1yoafVw+Qbo0QmLOVhbI99D/1ckJBKm5zJWVQ3/Z6lE55qffeIHkZwnL6LVJ3uZbsYi
KRefleZSrR0BKQ92fTS6VY3N+royKOe9+Dg5XTcZkQHGoTmoIkhY3umd2Zz8mkzKf6DwUrRbcn4w
wd5KcYNruiZhRGJAuZddHqEuNGS+FnkSdXtcIvCvvEA9yk75GtTUbDMHop2Wmv2xYwV6qJ5Ahu8/
wjL+s8CIPzsaeq9rRjIbqWEIyVbn05tbpL5NlXgPfN3dB0fDkkY06KLisATlADoeKuxeHoUJgXdN
BfSr0v/0jO6LSnLahEHXl7sQEfIKrUnm6/LeBs2d+Jn6zg8/wG4ZKdykz5ZE4YfKvcM0QzeVQuhY
PfsBZJz+nIOAwcv6JPre5UHnzpc5hhW6U5KKQnxN79Tp7ggOQ7zH5CkLc907sVUqHhDzvewAaEM1
tRox0yNdZKqUzCszPNPTJ2bJpPFLdx6DcugpmzMgdF7vySfQmY0KEBTftshKElF3T7jz3ViJbS/6
2OdrzOEXZqHUMkFunKC2A4FlUOAtYyu8KNmCwZva+Upa4Eq3NIzThZni9ijzV461R20MY2CvPAdR
jNqSiHhsVSXTscB8ij0hNj51oSnuIniUdFtzQcQmiEPAjJQ6YT08sFmaxE2kkGsLE4b+/mSugFJE
pWHJbtE4B8isfkrqChs3GE82/W3yGq1sQp1XT8WL3nbrcLSsr0hjUjrCQPP5N3gMx+x7Uq3VsmOG
+ptX+u7asl6tXMyhMBo9S1+nMMJ3sEG0A8D1aTbByPfVX9Hj1uRIlBCcaAeHC5CYZLHbCVRpFWCD
cHNsZZe+/7NqeQbHWnzMSK+6WyXNyDz8MUkssqgElBoGQO/V4MsgMLaJM+4yXTdNdHDmWW2ZyNZb
13WQwzEhUZ19Pba0+uoKQ7gh11eqRzc4NNZ/AKADdd48fRQBtaRmRqd2N78NOiL750+KnMZuz6vk
WGPeFHtAWElvgcG4XsJJ4dkrPodHUQYszgzIBz/IsO3sohEBV8AV9K4/M413prauRgbm4tizc0Ma
IBPobhoGUvrkWKR1KqZm+idxTDRMY8FiT3m11t38f338sNHNAZYhPUih57ICS6TuHUTFdq5DU0Hp
xPHlFCwxcyoPJ9NCihw+ZkSmmNbLJfuILqVRUH1yJndUPSvjPbw8kZG3m1L2wLaR/bft/xZZ2YgX
x4Hfg/u4XQF3zDSmkUaxkWGCzgqNmqqhunUDrvnQ5V9y1tfpBJjUZXY4SUvxTsyCUSbCzt8Dcfpl
47ju0+a4jCgkroPQupWXrOBTGmUMmehod+tx/+lG/dFejYtT0rayewOYGW+xQpwnUkXXZcN84uWc
rjSPUGKYgtHnUCbItoYwXiVgXInlAzQOICPpn44n5D8+aT3jNRELwl/wxa8aAuJjPsCmqHJ184Jy
Keo8civsPTqki/kFuCmk/H6TnDmh+5YdVbYmYF84oQWAOJ8dCUksxoAD4qmJfiQDY3bCovAl7YIi
wKe+FHpYaWwEA8QwACPkxr/oRcJ07f2i1tcEL04ZdAACFABP+l89orm4JxNtuQPykU/qU90tYvZH
G5073KDDtn5osSbyS2eNyQsNwHIWEOsn1lTB7gznQXKzO2v+MsBtaIPY4d1l1nSCAFG3+TF9M+xs
CiSG95gyzFeFhOwrhKNTry8EuX2ycmnzv7VqKO+c37e/AOLJ8CXuGkFrd2EYo53fNVcafirdqBDP
S5jn/v+1aZz8I88AC8J+yHwRvAjzrr9COlesDE2jxEMv5JTTsVi8NVf8UpiFDEx7NzOPj0kmlYUO
EutpToTqund+XHQN3T96iiqvvLUgupzW4G6egCE1EDGVbb0at5E/iGjrupcx3yA8Yn/ugtdY55O2
QOcO8wvsYbsxHvB/lCKzy3SJVPj3w7m2bbpfa8eSmf0wXxTEP8RHPF4v+UucEOCkr4kQoCBRY9Eh
BigjGl88c95yQp4OMwS6Hewm+OzB7RogN7rxXjNCmDZcfG1uVySz3ZYvUrSm4v8ie4+mM+hK3C2z
myWE+CKtAvn6vmPHf2P4YJ0uWo35K9Fa7D+RjI0Dz1rZDCUkzOpkZAl4Co6ovRaQdATZPlWVwUV0
8b0KlzNYERpxhpEbfOZJedseSYrb7c9EByRi3kY1v0nXxiIQObpLi+uFWN9dBvKf1QxKTO4z1x3x
Siro/LZiYhmStWqIq8Ks9HAtq5u+5pcLrhwQS7v8ZqImmpAjTXKdrkeOs30e0e22BItIIPEMjz86
jKl9HzMH3LADVo8yUpcVEZ8comlI2c2OuQ2nHdItIP2AlmFbaKRneezU3i8vEZd9yTQlZqx7tYoa
uedoqVasYDZPZYKYzDbmqvEYnkhLxaqXaX9YKHgw+e+cymwaDVJivLrOaliXPca7z0woIjC4rLH8
B2BCStgBaPCbxSmyZW9QZKjmDkeG9frEIWQd5h2/yuIIr9Cyia8BzqeThZWt0L01oorswChlMPfw
lmxXv737kO8avMjRd5xJsXe/QFFb1WwMqq4a9tTxHGQ6NwH+jgUZ35VTlEXYzG+gNGxhuuGW1dOs
rkaQzM67orkW+7pKpsCHJ7BebQljME7XiAuqFgowV+LYdKlCxArojQG1BWL2NWRD+6C2vnml7U+g
v2gUV97P+dpWL/2noQ/b0O4eKTea9XL++JsJ+mD8f00j+gPwrW0IrA9rYkJRh1qNvigxAhKkeTVZ
CBzCOY/MJc6xMKlh1M1Vv01i7ULeJDx+gwzRpiz5p4jMxCsooNzGZ9lAGYrTnoG7rNsAZUsKsUi7
lzXSRvtSclTYrSuNJqdYfyaGUlBjRjpy5yOK81cvE22hOopil420AtYzN2UWeNmXYeZw7a6r5WcA
e67bgHN5qVLr9CAo5ad7Bi3MpGXtBIcYXVVVqVJWgA35c1yIPL72Zqr0NBn3jptzRGozla2KVT8c
jvrx4R/dDdj6Vk14YvsUc7/WLZljyCcoDihYf0l5m6L6JRybbt2zYt1btk2TgKjEgLnkqjXHAHqp
xyGByk8tb2DvRcvp/23QTTbxAfaqZsatqG9bQuvsYpN/1uLT9Tl++pT4ss2F8awRlc3kJwnG2njD
37cNkci0PUE024iqxyTkwJwvDw7ANmBueeMyICB5tPTvG9urhqqlPKQhXolM7hn8wLb2VJVCZqJZ
i7bbzORcX8Rksc5MAxFOhoNzr72mZFdHZHZrHGJ7K+uGMLqKpJS6jWxpfUHGvekgJEZuApBhX+3s
NGVeRmWtuwwR/cKYQZrSmynXMl6KCV8kRMyu/ULJHZ0lLoCTCVqytoCmhFz37an54xnfv4G1CUp4
b334JBeuQf9kUVGZYXb+dzyKa0hdshH35jg6Gh9qdcMvS6/BYwlf1JIuoybuPqKad9jLulfQ7pFi
f67JiT8hckiREH/MXg1ZQ4/ws9pkQrcyhIi/z9jg9QB7hrqelFD1calhNw4OER5KNUpp/T58dJzg
7YVW8oGIGVygiC4mt2u/Kz4uYGtYYnp+dL99hIkjuPTeDC4CduKNdIoZwkm+cp6LpKXBwC/lUdAj
duSFLqTfb1biUpxQpQZlNj65YWXHcLGaKnOKdrlbLQjxvk7fFqXDsfIZacSfgfwKUk5r33yYvDPZ
GHGYM3COVbFRidgybg4wRvEy9/EJeG7BsKZZ1eSg2z9/zbl8o/u7E19ZvOi+RQ5ACosF5n50TSa5
kXXixPpoNPcoYiBOy7ureyLb720SMOq6TJST7neiR8mesaGoM6ZrBPiW48CbEUUneE9Kfn82/RSJ
ZYb5zoc4+64z7RtPigzwkafLUwg4lMtfB06jc2B6+40/MQTcEgNMeOYSckN3zKyiBtIkX5dHIu25
0L+KgNE5K1l0FmLpCBG/Zg5CADICAfmW+ytP4AKioDbyYSsJAwT4Lvx2i0rhunVWzVU1321ohy9p
stcQNfdTo1XjTyL0A1yog+5ay72xnqv+CV1NWqLgILbydZCVsbs9TL19fqPF3doq1Fv4DjJXn6zj
FvgKE7jEzetKB5qcBuJmwkUaF+6u+sAOn9N2sUZxNQMsfZSQ4gbxRbLOl7hDc+zAKiNl2SP4aHnw
xIpwAL+6RBrSixBG73GYXRCGGodM8MgbBq7WpLryBNk5FjlCnYRxzlTdtXK2P/mjBkZBZxoVjp1j
lHBKrMdm7K8N1BL5ClxffsZMFyGpcE0ZWBgvPhAeDgURU9qR9eQhn3Fp/vEpCHvYX5J0YXVqzQPD
4eVwkB49PyImAU1iSNKT7TTRk4deUsdaAokfYrg8682fzFv7Gwy65RXJn8gDs5xqPTsK5QkmSsy5
06uU37c7Oj3BZwIh7QAPI0dbxPXooS4fAmGt/l3LYqvg/OLXEm/ZklfZ5P1BdXlDpwG6PAGpayCf
3b19N8E/+9QYXgzgwO6Rf9uQIlleoKLMCVGuCOIzzmqc8Dw1XBM5+qsnx7tHCy6BCruqRisAMXYp
LvOtXE4fjbzRvmQ/EAuKXRGwFtl59g1HXJmE/QMcrSTBhcEn34KOSidVdF42RqrE7HRelBfPdk7T
Xvq95DhjCyYOc+rspHEvMcDHdogVyT0wTWY+SpcgWgAla+eE6MbSvDYqJfKACIM1WAt9nX/BJK4K
zxwtaS3D0y9wK8pDLqjYiiGqyXyNgN2isXU775AU/Si/y6892htQtrsLs8t4hu/Y7rS4IB+tFQoE
RdAJ9CGleqFhZWX9DdJWvyeMN0v3jrm4km9QuhQgRiyvsADCrVg/fZfWWN3aHucDOpFVTcPSWh5L
Ebd4j/lBazLRkYjVCM1GA77DbmA0mt7ATmhCwhNb0fR5HeHapXr3lkkNVAsmZSlM5ZMP8OAxNNkF
emC7sDLgbRZTDlhMUvBV4NHPkv5N/jdRlJoSPI7RjUefDv32Nvj5u+zeS5FUMwcoCJ3iMrOjSUbK
QfHoqOUqJLks7oALsCHUonIWL21NtL7mrPPAR6jKNDnIvzHZOyARQSSdnAXOdT1GqAWJadWm5WlI
XTXXJ7AkIsgutKpnZ3Q53YM0bTstuB9qRqzV5KtjgCqyQ4VZSOjJaR6HqsL4TwPi4h88ALVgsdqW
HhY/8SFGIPqzulD1NvLbU6gziD+h208SHufMwEtY/JcvdRhZlKUF8dKBHEI1VezCUtxHtXnA32xZ
EJvUS37wc4eHKAVXJgo82R8ZsBX9iywHzqEPLe9p/iFzc7QhTuKYwNmeaXa7TdvUZaPLFRfI9+69
1YgHA1P3jLfmcGL3KcyfOye8ZAthGM8zqrvY2TETMf4kEC8lD3DlQphIR7yM94NT2ADkLmphtl44
uuP7NMm1TEikefAyX88+J1/stYEJpTo7JhlJ8lXpH/oE3BLlbPYh6UcPv76VTlJj8y4GzFM5UX7G
pimDiJ9GQ6pGD4TqZDnJRXmEPt6qzhf0v6iP9IKQ22DFP8ZP+C5Wy9fgqn1xS8zfkLMdaI68iX8Q
2qdbl7q4F1VAWAV3teH+GyvrIP3qddBOBiwIbxDQNQfjlHKZt2nnO16bBjeiFZsV6s9Cwvp1DYtA
dASvCcL0ISfbpnHC3q96e30EucpsMlK8qiK3jr2wAfMLt0IlO4WXikUHntsNWNohZ1/YsD89VmWk
eRYMxzYoGVAvuTH0BciKquDeZGMQJKY9DmUE5WewyZAAiUlB1BHFKY4oM4OPiL+NRg6oqbSWYuZs
RsCuCcnHg+Ge9aEQ66VOpbtsKaFWIpupD1kkP85XzdULuT7/b/g8+i0qnj8eTBxwKOb6uhVUPnTs
4Vhm0igSktMeZnvl4yhqpBP8HtLhLm6yoNrlBnCAKEKtET89pZcwV4+iaxwhbJ7qhShjcD6ZmlIZ
bDV3QBsXo6wANTQ24EzDy5QNjBTxwnkQuMQOJ/BzrvEC74aquEY4cq+8l9hdlTmK7VvcEUFqsW08
WSGzN+LlMWDUsym85thwFiwXH+URGgDv9t6hXS91DoEA+rkBx122gY4pOWHJI3IFmL670det3XVG
iOzuLw/c1XtPVENm5eFV/JYr+PF0XuiGiyhJSdPpZsAIVS45EqrV2B7oOpUTkCboZRdj51SUAjEF
vFeYu1GhhspFxofipiweI9Zy4xCH6a+rpv+jSA9mTj0HURiNjJunrzIIR7Wq42D6aqtga+8PH3uk
dNWz5oBgAZgN0Jz9OIOsCYc6E/pbSUqWW0n2CihZ3B+PycSncKIM+KiII28ySa8dHkXkV2qN09fE
O16oCWpNSMEkPTk8bjvyTbE4YQ17L2OPrSJ5+/s4arw65rsbrXiMT7xuEAeaJPPkrjO4d7LT1Q6X
pOYkjdryzFjj3eN69w538QqmAqVnQDMVxZd/SxVCJz4BNIAJmgQUcStBN1d1IH1ZGIRba5BzpIRy
BCdbw0yQaktHgCBrAhKfS0iLhvYyl6tkXYGgu0grR3c4ZyQrdUNP2gLili4Cs8KQ4DTsFB5rDhpG
tmfmlkvFtFlgBDZOoZDV+mc7KEYjUEGkNqilCmrmEeSjzJZcPfi7Xf6zJ9SM4ubzCptz8bZ4bNyR
5tyXUALP7GHgWoSlTANBjH5pYjf73ZA96SWATkQqM6DX6SQVdjx/qbuRRtnfgGcuJgl87BvY0EE0
8NAj0Bxeg29RywknT3ee3xyI15PXGFfy6fVKlLCfgdC48PB9zfnwzv8iPBw2U4ZmiUILJfl+00F1
HateAI5Hjdo24riK5qey+wdpjxE8NA5bKdv/D6CQfa7uecqpNrk4jUlTcS9+b/+gK2v9jqynKrak
tIrVCVyC1BAAOopnnc69s4u47dCORECFztKv/OmKon3ngiNeZikx7A1FzfppAeQwvqXFEwXQ7B95
DVkv/q3Fk311WvUbBFw59+zJgONSDWmIqdYmZiSWfBZywnGl78QMhbxekgC8TNQdwDsetYGYmHX0
/1oOo2XKActuKxAg2+ihSzlrpKjnWNnTCqMtizbNFZoq8Ltlb7E/KPTP7Mgnybi3A6yFlmQFkC47
NXwy9FlRJV4ooSRP3jL8SUFgdh9QdvIlMJz/Cv3UJb3B2ttc/LzWjmj1qeV/dqCpGg63cw8AM3e2
IGM+sd1zDPOEN6C2ZQ731HYu1VWuAzUFECF6cr+1ew9Q3BIQ0VHVOc4GiqygUErYhNSExgRFhs63
AnBIPpXlw/i65QtsFDAPJoWQM67o7+dcjPBIKyr5/6HNRgxItxmFvtj5cIVF008kD9kUWErYWiLk
mPjd+xpvX9odIwEhqp8VspqwzfNSLETEqeOufSL5UdOzE37oUzEDr3ytS92SqIQjL9ejoqhALNQ2
46N+zxGPlUCN3XKuGg20/dtgb+OOKUq5lVN46m/7QNpHI1FbBw4s5W72K9/CKpOLiw9QOaLBdWWF
9CGw7+x3nyws6/sQIkiNQZKLV2bLWu3ExFv2c+e87yI0IQ16BAE3oY3RnjNOaAgOrZfpLcwcGvUh
g+rZBF6CeN42OOGR4uPJWEjH2Fjv1BnRrfPTxdTmm4Pu7Pm18J4Xy+hDpsTREqvMLCr5HDiPVb8C
kE4dM6gWZBl+4bEHv0q2TKugN7Fj/Smz1le03iigCpHn4vrpC+YyPJRQa6va8XV3CRo+76QnrHQd
4U0Hrz4v2Y4gYKJTxcjtVf4zxS2JNJEV2nQZ3zq4wrwt3wu5jPW9vluTenkrXGteH61ASQ93qt8j
lhyfdsYFlYZFNwpcAkBlagpbfmjZp+5gca7WSgocvSi+eB6SL01dFiRaOuwzZfeu1QkiwB6KvTnI
IGX6m0fzhdDSNR0ZPJWoJdMHtb29GR5MphcYS43iXK+7dCubPTMzEGCDlH4UZCkAElTg62AIH5/k
VrmVpZ4+nboCsZBSf+E/qj65eFBiixaPjbkV2FULw6krdAEr39mTTQ7wl8IOqet0+rVJ9pmvdrJs
ZpuuSNC0Ss9m3SnWfi2CojAQbeeXSnfj7NE+ZoiAbqBjls0et68TfqPYjKmDV7FLEGumWV0LBSEb
YGw0nSvtogcQQJN6nzMU2acmmRZ6gV6K7ldVUqq7SoedZDucW2stSHQxWZgPQOauvHlAzLocj2SO
4dSRvgCN4RzA2RgWzOykprVBzIuNO7h+HARRrICkrU0eHa3k+NYq1I9gUP/Owkjw1Hfe0+vu7bvA
mWXyyozybb3+gUYQlNOxkB+Ka1slzSjRI0O0MIRYmABbh7khD/Wh1DCHsR8T9gR2AMp2VquTteSQ
BTLbmZ47br1Wf1iQGnPFxPKnuSYljBAMNKE9W2dwbIrRR5Lya82Wx8SDDPPxKdD84QooyGqzv0re
k92LLjZ9DbA7pPxbVqicY+z16wrIpD6P1h4oEZYnFHwM7HHfQ3Wr7YYeSk16PuBGiiyYSRyHt2IN
7jVaHFNNAfzP9gDSyq5K/qmyS8yO7e9C+mJQTRTh68F7m0eR87IV+K4Cuwbp5f5cBfiCYHfXm9I6
rOL/aBjCUveVo8dySdAw1NKeN0X9UzdFmjgaS2qQApv/rhIUPpqwNwLbgrtUgjwR8bblmhWoAeTd
E+X6weQ06KPQMPoqY1ep5a2YKPSj+IRobk68n47rq8t/Ay9lRsENGXxQccgPtmituyNYqmfW6lSI
JoImU/ML5ZTAMxmdINyMY8tCo+7nLVwVTOPBji71mR2v1t/ymGu7uhu+/j8+k1rcbbPbD3fcb6x6
7bQFg51trGzbj2HoPhnC72Wkn8ZQouPZAsbk/vMNkrb5WDRRnFHOD2TjvvmzfgnpgvBK5ApC5/WL
vKpjGOR5QHuDDl8I8QbRErFdRXN9BiHjHEojQwXe5pPkghirD2w4+lDJSmZmOfdfRh7UQKaDaOP1
5H1QM8AJhVvFyXnRQeky66ojkMV3v1qzsVTP4901tjH+2UOZpsi5sbboO5snq4rhULf+//WV28bk
EjcqvoddjDxKpivCXjF8H+9Wlsz4unlul6v8xjcLMR8NgBChkcK/JHRG8BBvmYUSpSlIq1NRrwKH
95Zrl+xV5BmOeF+9QI2VbglFbuD0Yx1xtfT4QBjAK/aVxuOyLRCR+zAWwZmT43eISz5jktJeEJCM
rb9eTxSY0jegZm4GCxIWLUz8+jsa9u9clCIuGUUv/Af87pR38kuy7Sk+69TabNtFSQ49wqiXGMMK
l/y1fCqoNqEiOY9sfzHQPyVxtmkLpfGojHK+J6BF9Wgk6AbMO7Q2r3Ls2vxwqlvznd2u8km/1qZi
3DrYYOiikhvI8vszVh/+D/5rKv6VsBsqttRSYOuOP/2MeY1/NNV3vQa84BtR3WEBgiPjTuOUOa+I
eNuaFscDgJn7+uE989xN0Q62z6KCKx0h9CScriMHxfGiIAJcxkqUajqAlYFCz+9lGl/YULZExoud
Z7Z1JPDzZ7/DverWzAI4fBS8LGN6zKfM4DSbOH34rZl4V9DZVY4U93ECsEHe9HYVG5E6q3tuIiMz
fAg75Qrkxo+xy0qHLzlYQlDWJtBu0GWuStfHVNSvRUGI7rSEOlr4wlm5IhBrNieODCKpJWA+FuV0
XZCYfAPTJGeyWZYHSgPEwYgl9otf6eUxsF8j+7hEOS0kpXc9zEACr6r82Jp//F2ec5h4Qk43mngb
DyNIQreMuvkYbS6/IKPQzr5b7EkZYR3bYIZNNZRe4cZgRLnbNPRT7YiJ1uA7CjKPJdDhLDucslb7
RR29C0bGj7FUDEDWZS01xikQWMGatu7Y4lTgG+McI+rtFXXQsbbd2dPglUqbGJeARBEJLDH2F9bO
qgZbSZ124E5u8xYqmXN0rqiNaLQ1qj7bRhuYIFAD9rtpZSpTIzOPnzTq9VeMMhfhrvh+En6JnGv0
PE8zP4UfylUeZBea8tOK4yiJ8eV3n42iTqtPoYD6REchykVmngApk84UnudZ7/F21xlQcF33u/ia
eUxu1mRCobmaaoiSc7ftbO7GF4lXHJ4WalRF7zWoOx7e1UTczAHnA8hmK/CQh3Vu7chyQtEnvmeM
+uQqvmnqRgxDOmLnJgZNduX8gOuhydVv0WtCTjFXuBRqquCusM1P6CYd3POePpFfdESHcxZIYN0f
7lUGvhxV7lQd1ypnqceu+ckldf1eoyHf1RvdwEP2HirNYcfPIO3tbeOeIwj06u7tHs2pxHp6AWxY
hVxss62G1xath+usArumO2Y4fM2Oh+d66WBRzMcZQWbqL4hGREPL6BZFTp6t7ErpKDngimacdhDH
KVHJO2tr+b5TDLv2XltGi4gg9SLaJivU4cw0dPRIRzmu+Q2/4NHOXkJpBzsJ2w6jM28lVR9s0wG1
PMIfSwxV7I/c3yGMNcV+QFiEnz7ccIiXVW7L5FiQzS52yGioDtDozT6heoTsCw1cnYyeYFZzjwd6
qzi08DZPiSZLsW0JjlncJhXh7t9gfJIcyqFuiQ6Gi/clD2bgjPYgjBUUhguitzOAM4qnVF2NgyK7
LjlHKNTtzWP6OhO3RnjKgKn40bVmZ9yeSDGuy/bpnLikPvbxePFIPQCWnfNPfHH7/zaqcbzmcq43
doBMKcz8xhsMlYQLjn/eEOtjNMELygiYdvjrEVlAEeVohobX8EfYpZHYBHY5WPt3f5eXaAMBePmG
jtkXRL2hpwKzmFZtSva1yOjtnt8Y4qrHplNPpgE+WB9EwRuGXa5y2dBu1Mfhg97AZ+KBNsM83XM3
SGdWegyJaF8uHNBIGpfPKW3D97hG1svh5/5T87cIydA+U80CKA5tokwkX+G+8PsCOr8xN2FmFAiI
pxrntrPsmTcJy9Ksim6kAijB/MBb/PhPN+h2Pz9/sE07xXaxZVse2GmNL7iYRjQReYWd/ZkV5yxt
7FuveM+8UpC0fjCWoi94yTepoGm/PY8/ZGtqU+crXMcO9dxq7/3QYgPIMD4U29yyhl/o3JBJtgkD
/HVx6WWPwR0rwLPzI0zEJvjQbWRXOD/FOZc3ztIzqIry6TSFMi/jt+ZXv4MYCH5QhmVIqVz1WfgN
fThuniitSwQDuJm/9PyekdN7Ze9T6oPR+tVA2sRNLCY+1iewcyou04vGxNJ2jjlTHq+tavZjcUgh
B228tYLS+lFCAzc7JVfTb1fG04ZsP8C73mPNTbC7O9evIsVL7DCXCsgPTgo+UEMRnyUGMPEyOfA2
07UqLFuBJKdw2+n1vn2QfnjG/UvNcEVmlEqnzX+/WJI89ljQbMR6OPVYMeOWnnHxuURv5thfu2Aj
osNeGEU70+C3F2MoKLkJOQaEWILsVXJpQjrh4RRHcc/Cw82hag9JTB2ZzTWAdKmfJ+jOGkx9CTiw
FvFomRWh3ohMzr/ZOPHpirlUGhQfAuF4hqzbRlZaAG5vvWfUzo2gBr4vowoEj7wi8hYSP/sUb3na
hrkJWGFAaIqKyfJISBkFibM7ezscKStBlFO1EIQkdpviFNQjQ98yNT39rCpNPDLHxvjJkrOKKx5N
AA5QQM0NVVJe8BalhqF6koHtd+khWwOATnWxdR6K1eUetJTk/P4/CM7/snTRnWPB3Qvw4Y9R6dqn
H0Bw/6WrObTVhEC7KKIckYXSJwFbhKoeSLq1EIkcMDoOJS9/97nV4QiKNbiwo6Wk2LIaHv6VfEiZ
r902MmshZ25zligzNnDMH3JOJRT89ItfPekoF/AMmogxH19zCQX0+nxzi5KbqdN38O2oMJN0u/9I
SXyBNe+pL26AoQj3g8d7BxmirbN5E+dXn6yyTgt6cqseguUIkahQ97Z6SOqHgo0Ppoj55qaBJd0k
W6b3q8Wlr2wsb8rJfTg2zmo7ir/8tPjgI9hA5VgT8jfjG0/WwACbn7RkuDoozSvNElxVRRySWVng
evR/fKwbyfb8nN9hN0fYbC739MIb2ivvR0KHwiMzw1R9Riid3M8ooH1NwCPaPmOAlm6Rfk6x+RVA
se7zXhB0FTmBq4NnrZLYFwAUdYp7GBhO5XSQioKuXzokqvKS6W5DTfl7CfROe0d17mtQvliQPWM/
w9VLCd+1uNbYa09t0PNBzs89CL7XpGqlVvQj1H451w91UX7uKc1HlVPR9VM6W7TAwA9kCXlJJpq4
8KxlVEZaosOzkqTAtdV5NTcRQoopNDsZoEORXuj2rpdTtqjW+4HPgBu3x2tfadXgLzj7hCHst+z6
oBzryb+/KvG5tbO0FReNW3g7Fc3sBLe4kf762gP6llenED8xeS8dMZFmfmxZ1FZ72ySGQvEWukyg
rMrt7g4gWJD7vM4K10oHmptXYxExxcFDJbMFdv2wHApNC/k2cJNSSnJ+93dROfSoCyDT4gUINpvw
8TILS3u36KmTY7NTgnVBqKfzufmeKyI1VbuRvnag+S/js25js0zBQFzcqAaU2+CI0kLSuIRXCbiq
NlhVjRZLLP8r7w3ET6iLvjLi2gEdEnJNktsRNtUJkshPFjuIrq0D6kQ3jdhXOckgV8Dry4bIyPXK
5rUBq9avkRAuZe9jpxk+JtI1J+TNonhGYHvVcLYPq+la5ZaWl9UN6j/TnwcWXj8Pe8kPeLPsmqtN
CVxZrA21kRKLMoE1m9FRSZhyQcEoMkGagL0U/IlrBocksoBfepFP3Cl8CU6RwLaWhgQ3oUDqQ/dR
OyamI+MdGwOeTjpJjpXYjjsUyu5+8SUEdHzafhnZwzeyHy50M3RdeG5kCjBPX8M349LRX6+iWw2U
GtK3LyEEsq0ZmP5RVvrWA3EjRUx6EssXdL8Ys/34ybS9eNIrxG2SuI5NSEy7pwmYx1k7WvnXsNnJ
ZQw9ObtBW55NG9qlcMUI5TNM2J0eUCpPTM+be38M595POh+cW4b7fEdaaMdOKRkN/tCnpba+DKno
l0MXo4vhTQQuPXoczLFV60VyyAVjL8AOvX21CIWxAlgDtWFECiXUaIPje8Oaz9MDrcBs0E9ns9TT
dBpZljSxMFthuoGzzfTQAa7NWQ0jmnblN90w8vV27JiFNb1eMH34k2GfxPCwA0v44ORxURbXhnzq
Ko9VooUI5mlLwvoebL63punLx4g1dCUmvWkN4RTd/k0K1O1e34vRhQjDFwyq6n3T3g1GAIhqboZ/
BbGQ8Xt8uWqIiQde1xWM9FYsua4M2p+P8rMjnaj6eOue97TI6NeDVZ/6d86Ty3AcMSBQMBTXMTzu
ie9YORN2W0ABLVtKnP0klzRqbhWupd4kCXX2hsWmQr6ASAXx1c4l4fcE/XgSZeWnTasOUDelF7ut
qH2OY0tPZ9n8I0k7Oz72tXIFaYej0TOhA+iQqttCifoyZR4IgpYvZjBFgqSqUBIVWIwHeDpQn9XG
0wPegAtFL3cqr/7IWEP9IcLg14gwX1wgM9HxkkaHputfxqOnu6YTjFKywRz4VqedWFDv9DzuzF4v
G2mstetbD8NKmcKVeBn7cNZOQWtJ1gvm/f8rTjDoev3mgWl/dxfLvLp/BSU8Nki76bTnXOyzPVpA
tlBi+wBqzSaeYShb3x/8z1I3I6SXre4YEYOi/e1Is6Utp/05QtG8+YL2lZIkNkPrXh3kJwXYeuQS
kzrDqjpJYFpDacVg9PoyoAVjTwJa2CVri0ll3i9prdV/0qKS264OGVRPYSLE9uJNIAclr6ZhvppH
TQTpLykoRj/OXyrooPWie8rhJM11GArWI6bUDlcgrM/8XMF9MPqonsDkn2sk+aKVi34ZyAEdslnv
7QyZ4tGlEsh7EQpwhv5tTwqnTZn8VFOyIkkVleU/B/OnbVPrB9j4MvXbzDw3XkjDsgy6Vv6V1R4m
mbVX+CT/zogUeqH6JE+Mmo/1NCVbZ9u7W2Utx24WuQ4m6F85evquUw3b/tp3Bfllih5rD/QeqzU+
4c1Sk36SWvabTFOsKhZGXe/REJ9+lJNs/zL30nMnx1rJhTgce8g/asf2zwzBXf7sOB2HY1XIY6bD
bPubRVIKPsAmQTrfRQ4GnakQ9r3iMcxPWpch3+M9uqRwmgGINByvDLOxS++HNfQ/dWg5/01fg0ho
OxjbjfrBYqpGUtcRAbzF7tgBQrFQY5UzotMbFIY+Yef1n1hGpQ8u2BH823L7S3aYnUZOEYdURyRo
69MdhrqvMGYbSCuuexUjOSN8MgwbmQ3MtQN5xgUQX8v1j+YDFpr9IEXEAgdbixEOVY+IkdQxHg7h
/FPFPe0n3J03/4Df27ObQ3jYpiNjqB1+oHK5OmUUzAYAL5cDmNYio5xavnIX+z2/7Ybmm/ZwNGho
XnnS4VRpvy5CIcojojignx1n8d817nVKpEFpi/MBHAIiHW8vUGUAjizeIGqI3EBEt20FTYKdsbfR
stASukodsIf2M1RxTy1GCag520HdaRACODgs8GFDoGRWFdT70Ez/VrtMvORJ6wOrK1RWD5BDCFZS
u7WjuG6ez2yACLIMZbYOA6CyVpZVyhyb1g795BcZlFLv3wL79FkrZ4riE6Mb7evPhXbSE5d4KmT+
NP2Iu1gVRA486hFlY98ILm1JAIjlEm+lQ+2YE1KQ+Joj6J+CFzXUeXNRkzKcWWZDgw5Hs7ZeuqXC
IyKb34rq6hhRD2Gr5JOKrqp43st1+0v0X3LRJnF//y5MTItKtAzGQKMYy5PtI65MiOAR5GCRQzS1
RTVjisl3695x0VJF10O4DSJhhaFD92rlCiq4JKELejxRo3LknyFLiF9yxPNHA5eKJJRoL7ktbdCR
VYyXkyGzt4VnRz0QJDUNmSxxhfD6FWm1CCQvkCp9YADK9JWdhnk9/piLiMLQm/UeBGvtMfOE1IZD
OiuL96QTyqpmRTUYvM8qfe5RSC2GDPo3RLNEgdxJBsqvbNVT9AQxKVZqgKLz4+7rQpUCrzQpu54x
JxpAkfjggD4ggbC7xPu4cZaI1KBiVkH9TbFWTuKW2vfO6W23jZ5ej5lEryEbMDjLVPTsqOwWNree
kKSx0MtiW25Chd7Xm9pZ6e5IWWBkYkPuakoYxLVjIm+bQ9UG3NwIofwNzOf1eaKUkLf+CznzNcT8
8T6hAAV89j96lqVdjkR4EuTO7DBCzQciQj8VMR6jzsWvx9QxVQiFSzY4/92/nJWfMcSZGOsUTOBW
IDNJ/9yZMJvMX4oeJGXd3L/UClb/kG7wVzxXw8O7I2/l/Kxe9m4dKC/VDAbicNRsdGXUK3objzIC
PSQbSGkAydJOwyZcPG0WQVdClApIUVK3gv8erKtwn9QiZtUqtgN70zBIIsukqVFFm5gIMfVYSEPO
oNgoN+d6AaUaFG+uqeiI5VsyJzcIwJgQSl4hlDux0pUOyUT33NMkDe7OEI6XQMW16NX2XfSx/llk
avlrflDrtrZfczNxahiGie0SPb8HkKtIW9Qqgm0wUivM0EwMYNfEEuMfOx78aTVXf3cpSMmNTGs1
OGXZSBsysC3AZmfA1q1ygqTlqCPl+StrpuR7ShASdQj3v6zoToJhX+TSJ50GL/MtzIfMWxZqndiC
WsDZyT0+Pl2z/FARTk7a0AuXfNTu4KI5GxVJJxx1on5UQLZOyKh+u0fhT8ZLQ/VM3i/O+WFGVGnv
F8iPIw1YoNC35hiyuK/Ih6wVbAsHSBGDHBqOpnqqDsAuHYomX88e5DVb9jwF0ypznDii+lhkN2QG
eCmEA/DgIf6frvTp7cYsV25rE2dpIaxZvajdUlMoJFqBJN94Le/UvPp3cO3sAsVtcB0lRle4G/ar
oMi7+D0nVQcrZS0UfONdVG1XVwGptxzLdiakMHXMMYZzhFxwHgXp926F5MZlFl94r8GxsDIJbfpv
mI79h+5AM97tHufxYtyKDxgxgj+rm2HztOOPCrtxW/HMbm/oGBGeYNwjAZKxxWXhxUwuwiqY3bxx
bYkWAKi7fn4u+EYr+DWt5vh7zm/DDHOtnKb9GPIwGa0pG3zAnqDDQRpuNiSBuLDjQTAgrs4H3RPo
V5qOiFGLuVFaOXx4JfUMD0pKGlMyqxnpcAX89X2GAN6lqLXh4QCKyjlmbZMmhjVrtzMXp92x91YF
dQgBEFbN9/5xhX+RQ3BFovsJSU9hj6rYFPgX/U75gDA14naABUdThWTHbSYxnTkVLP1BmgGs3tZd
r9GbtaRyxKrlGddwEq/2H6K/txtLuOf1CpGHJC/flwuKvnpH1px2quuUVyDq6u+g2BIrpnpELLIM
H1YqNkwyrumPhea+qmJmo5kUp57Inlf1M+I8HVP1tEatDoAZLq3AnQBz8dDIvwTWXs/zr7nJzVBr
R09+3SNZSDomcJCl96tVZqOwoppLAArKCzoYVhG9KcbOJ/2NwqgMTozPf6frVEU5rAUo52Cw4aZN
b2+zFANNouDPri6Zjcik5ziWB3tWCTSvT3iHL22EQLPTj7kJOG7JT3+NTGmDCKoLielae7Xdxsas
V/yRsVYsv2Yk5bNyGO2SVWFhoR3lJsB44dlzha3jSJz9ghq1NPOMfCIIARsqTPDGxh6ika1R2eB2
bpqnFpllZgNFtPAx05EtH3qPpwZx/nvTzso9z5/nMvFHoWB1mlFPfa/maON4MT8/gEDgYVMExTT9
R8Lxs80GwzkbngOvcNV7RjkMbZgbeUYAk54onZhf+NPx+l4JOQTyk9bp6TjzPwogMyIblr1hDvUo
Ko+ZhIcpK2hgQ7jqH4jitzcYFIdeMv6psV7onLIjntpoRYzj0y34jgVsqoF+DulWFnFx8hv4tTMP
aMr5hAnMDDVzn3X4nMFlwXOJTUAFf9ul/jHif7rUqDFcvHX4a+qAwXoFMhe/8Cand7muw555rGWW
OyIyDVLOxbjheI9Fwex+njWZfRQ5blEblYciJkW9S4mrhMuRZHrwcLyNEEHa/M+gCmdvS3WdWna+
EAMx2HJBuFhAKcvEEScZOgHrHn1oh3jmjjER5ToPuvWJ5Z4SuNVX8RQY2cEvSDbiGSUKMFDYGUgY
oQb1X3ZqxP5xd5ZV4CgZpgjKLHhLU835Gd1qF+2I24jo98TpVaxcJFJlNXVOJqTelXj/nUtGdGdH
NpPhtKrCOp7Mbd1W9C9rkI/i6iD9hm93rlqgHs/m6dwm5PQ87oSKfuiZYBE3ZUT7HLuWxN/4+pju
jCXOK+XHEeHOjw2lDdZIYSdiViXDM7MMjZN9bRqnQpbwsTnwWOs7OqPL51SVv8ZgxYCwkjAAqnb+
tq1+QRsB+NYgbQHClhnPVJMe+6zBeQljMrQxrvoOMfIImBXLTgk0g5PAk363TukXhqRse2m9V2PR
l23h3h4mZrK6ABddPxCkL4oUr9JwKFRrG75ojzJqiHIyxolsozRI8zYiCM5HSm1aH/G2Ph7JP6nx
RDqvBENbuhKVxjAo2/bzKglG85mAaGXy1x+UuPjZFxQllspHT21DYAevVVycEyh16kcC9rHXq8ok
jlPpUJyGofDYgGGyU4BHo6fFo67BAD/maTlXpLgfwgEFZSr+09XAqfIhUy8gyRFOjZiI2vF8l5Hq
GtFN3FXoHU/TAeKrwcHYn6zmCrLKpd8k+ICi5wme3VUCJF/+v9dmLk8/JiNnK8L+kWpJ7ODJbgH4
ANXNuhkZLmoFk8/lJZBHeFTdLSiYvPI3yHM3VKXUWa2aTkAQn/sjBwSyKmHEm94S2BL/cIID1b1e
CZbnuLET0+yUB8DKGSEyD5B52rHh3hifGntMe2pN9ciFon/vPuqUHP4TQR5S2UxTokCyr6/3/Wk9
HqtOfNOdVIs0ycU9npNp9IUzZnuYg88KQziMMpvsiRZ4buO5aE+Z/E6UK4fN7bu1/rr3lYMLw4gN
SMuo9Qcq/nvKN3+TvVzIS9vO7ze4RGQmWp0O2qgAXQ1s6T9y5JXPuAGXk389SApObQfp3A5sTRpy
pptA7s87JURn+Gi5915t54YoDWIuJGLr9smT0j6vAr+v+RiAMmd9eZpqffwJCjvWCXLQGCLoHnoa
yyob/XdBiA4VecmSmEA+aTKQLhpvDlmKQZHhuPR7aMFDKsrSjCWNsnqqrCRXRrE1u2dXN/ByrSxs
q7qEjp69djm9lqzcijiWvm6gZC/nKPLCNsNgIhqWrbAqAuomQj8cl1jO1TEnqMTAt7H1gaTR6J3q
EWYYQqlrTOd2TQDt5LrNs6jH7EkapR3dHVdZUIkaaXXhNRt6JcbFityEfw82oY9Pzd5Uy5vN4bBV
tRjAutO9G+t4NZcluin5HGlS0yD+0yX/AV4bMDvh/7JJp+V5w84WE4ReIF3VT4le8smEYL9e3X89
lHBSuJ10s6JQxEbTsZFnrQhZ/A8hk7kt4yvzMOsjJDfIErzTvuswweJnojxAP7jfXk8fGKkqJDQT
ZTyCG4OcIj9UKOJakQYt4E7Mt7WqgBiAVXKWveoI5yF/xJv8qSuXA6ND+bpm4Fvn3VyEEVY1KD0G
5M/mufRnCCOpVfIXjExWi3MwdQgwWQXKlXLWod+2Q1U5N5uwzpFQ0qBi3/y33jNUIqkZ1SqSpdWP
gOW2gAvbDKdjBeXhHLYlnER/RPlqe6g+ieyc1Urzyl4wSYQOoARwbQNGZ3wJH58UfnJeQdedNUII
zkLUFtiEPDq3ksml3Nr/AtlXuoZtXdm06Ib3XgFNOKbx4tEWYZMiK+1gzigZlIsa8NqoQQQqREwp
wZAxzUQWqfBljJQHoURyAPEAYD9PBGPDWUXz/yfTbHAG0Ut5f6f77GT5rsn3JVZHsECYZgCgUFl9
kAbV/jakfNqM8VXZgEgo3dJ+122KC7CR01mUhRHFx9WB0ceVA3Nox/L6LZ0nIPBw7Y8124I9eZtM
YHGrR3pxxgbt/KPAiG2AsUhVO7RbETKPrF6AJS20z53bic7lex8DCI9keqLURsGcSe28qOa32iv0
qP1B5pvKYZzcncV/CNKCpMo4ZD3J51RoQxJYtwyNYG8R9UvfjLtz+BGeHNHxfNp9LsZCIhZptn6A
ByHXxLT5GHJWVwqDhKKiYBaowPJfU7wNZQmZebgXOmXM8h0gU1D16bSKR/Hvd9zmJEE99ZIgnkHg
3AhlKUM2CePg+15gKsvVf894YhAPXag/eptIIzhiTJkPhw4lTcTFc5EuAs0Tfg56Zyvl+FsbFXAo
F5FmN0ZESU5hdqb706+FBQ+JEjZ7FlaAKYcjIGQJMkRD9I9OKPNNDMdNoWCZwpb6A+IMKgi9hAan
g4nYLXeswjx34F8Wsv74EgSt4E+ZEnj9dPB8+/tgoPEJx0YW/L0cSEPElreSWo8Fi8edM8/evTyT
uLIBoWE+P0/qbPs8ygFapCGT7TVY+vpQpGbyOzFoTTDIaqXW6r5T2KHh1u5wz31TntSqrH23Algo
andz6pDwOyUEw9bG5YZVmwIyd3ruZWs9tGBBPInnCQo2AcFTjnrkarv+oTRti4mc3PSlHxXfq6kT
fVmcptICoB3ZG0YUFzh1f6uaSC+bo7MgNA60ZbHfYPsiL87w6V/EeW2kehrGfYM5yDFjcTqrQ2x+
Vin7egf+zzK8BhO5cL/PbnqNqB6RPdfIFw2YzscRYCGZejxawbnufA44pQVxmYCr7BN+r7KLVdOs
4VA6uFqbB0U12qbP0anJuhAoLt1CHFzu6P0OCoaV5JIMFNVVT1ny5Jd3XGCLSKLcCBXGOZRXgL6h
EjBtaZl1hHImNBvvgiEBYMbWK5m9uEPwqufyKoz8h7As3jgQ0tJ105uwVA4h2DxMcyJOXnHeQ1Yn
Fxx3U7gHoeQ0jZcdwE2r2O4OlcNOI7qclmsVSeBAvpacMRALasvp38jOurMk16olBksmbsNYM2+2
a+2L1oV96Ze0AycRYYX/vm+Qs+UXbLDvp7bLDBDDbJeCCgWURktdSFcxTs4c4YVvCOKyKJRFm0kM
9aN05gXJnUkJ5daFeC90l296pwMey24x1S6oQXlJY6hukdbhwPKQOUiqFQSfLfBD5Ydwfj8pz3eW
WDu0oEIsvLGomHn2q2Vba94CiWihkd7Et+TTg97TmLFX9M9g8gpzep4c20MPz73VgVOQ/6jmjIjd
hSVl8CpbISADq2LlnQjV+9vEAUVY2m5javcl5R7wCqezH2Km4G1cFWpsogEpzxVzu12Ht3NEL3Iw
PtJeHreUoBC5DTV1sINOtDnDOd/yINkfLPFZuvho28XECzwB2qy+c1u51Y/Jq9QbgFCPcBlDq0/H
QjppTTtTcOvJyV6BzR2eu5Nl8kf5qe4xoyybUKlj93RwjXM/mAz+TwXthrDD1yMbzh1ff3150zMQ
HmB7hx77hmHBqQhhvV2OADZFWkjG8uedso2+Z1utkAwh05l82kdPGMzGpnvMGmwhzad8ehLyEL17
UpkL/woDqM1IbuGqIjO1DLEoCdwE+uqfykXXugrmz9FG673ZQbD1IIS5m21y6PF75ajmUoeHH1l/
+3/ZYZegszM3celZqkoMTKJsQ0luXt6DOgqMynj4AD0eqviOQmpD5pbkI/knaiR3jNiNiyUIkyew
j5YEwVOiPgg8AFW+iA5QVYTbcl4EDOwBeBDwpaefW4UFFB820RgBTlO5PQlChfz2EVALdq+IYQ/j
9vUBA+urGfPIv/cr6GCG68anogXCd1KduJHQF2yoGlNlUa9IPLs+FOuutlDWL+sCTmWHXTI4LwLi
L2Vz5EujyfVoyXJTao4Eda8d9KUSY5gz4PNyACqkIG0dsh/EtcC+YC5SL2pTATpWVys9bvRBHHNa
UuU9hVPEqRbzgygh+gIr8Cbtbl0HntWjqXgFrExPs3TNo1KHpM7nFu0ivzdPb3EGmDP/f1kFLvTz
ovsiAqDMU35+V2OC/GTBCaR3eO6T0waEvBj80OIchFs2HFMpg+MgPtCbF8nUCUqk3MVPTr6+OGXS
SORMHRjWy8sZkeLpIQOXI573QIvS4wCm8XpdtWJ/Shn2qIoVZEG39+DuqC9WGHrwOZJZUBpdhJ7D
9gNCrRMM0cHg0/5WVtZGK71rs5yG0/vpjgEgnkbGV9p+iANo14HdSxo9S/bI43AgnilgV6yT9ygM
/da4TPEfr0nI0fZ1SUVvG0JtrvOvxtNOFNEZh5f1k5JHl97lzHpsXfEFjU3nrgcRJJv7A1MTr5c8
0DlcYAJdLqC8XaifuadnVQjTCzi+2QwA0+EvftaUQSLdFABkflFWp42awNs2hlRFtQXZpP0rcC4f
RRxv1yHHmQpX2biMHoA78gOOFDlUS2PM4yygmZshGPZCnlgCtYo97stT0mis+8fVHAfY6w4Gh2o8
80XuGzjRZTc+7759yV819AocOpvY4ks52xXt3HuXBdyrUno05mr0uerNpx/wfKW2ykkV2AJHXErC
o00yhLBO8ykm8nhiNh8yTAhCmLKE9W4b/AyRaG2zI2myQ6RQdn8Ry9ToS+LuYSFqwlSirnurfMUr
PXgImbVzNlv9Swx9f/3ucuNqLIIXstKT1M7EM/wuQY+Uk8c/mZq0se4SjUHqtxDI+9p8edceSCjP
ymt2ElnU1K11p0m91KHM9XJBpgZkQUmiGhMDwg5vFg1DmNKDwr/oQFuOD+ELnAfKWfBJVnCH2HsV
HaUA4F4CUZUnMIPfYC5UgboOwPluiPd96Pnp1krnxYCssDmphOWgTBYlzE7Pb0OOsY4EOZT2h0Vw
ePgX0jrCTSNqd+nRlc09tpRwGXOar/AMJLBvld9QaHXo/iyhYR+8hasBDYno0RSNQbWdk4bz8uoL
dpuNP+don3qeooaBJ7IYDOFoFivi6uhTR8zxP9FCjhl8wS3Sv9eqg2JJX8eW1gPfplT/zFPpJm/c
2JenjYtqZwLctA379ncl+a/q+ibTTCquWmDxiW5kSue12GpoOOZEzNFFKVYMZQVSZbVkoZLPpyGA
9/9doHt8QZr/4T+sEm2jdMU0D7uZpEdYwpaSJqMxFcROYXi6hpxSB7QKsKSvj2jHCWrCQwgZa9H4
6KpdVkJ732QU3gCLkSPHNOf17dyrKF4mOX3xLSCKxYRC1zgIvXyJ1aSZpzvKt9+5wYZf28dDwboT
pijrv8v8kzpln2R3MtL+sF0gti9YO3ZSOfx8oych7RIu2dJzplb6idDnTrrBGK6sSDeSsmPqok/m
44T0p7tXleWpz9qdiYjifGnQ/SDZh3ZRPMFhAov5WZyxFnCLpSAada+CY1wqSwN9XdGMfJ5G8DY4
hPNssBGJuAXCRXB/EZNNWcsmkmCaAO4m1C5g+4UQpIoa7fVlLyXOQIYmDHkanzw2FVJ+g2CJllnG
vaDxPCrCo6MEXWam0ju2/pkWGsDJgzE9hZfsVHinFkLtAXvXF0OsQfcFzyy4pJ4mabVXA9mRYY2y
VhtFe2Z0ZSte3COC6T2WPNFf4FmiyNo5C2vh6zfj19AkMe9UePe+l7nzG8OKz7PFPeV01WBnEgDo
EtI4rNdXxGxa873nQBNEHmSUQErFqp/r3Hb0NqYmWT+28SjctG2zsCeE7rrvvbO7TEobYfxgZmrZ
DITVrHSJCOwbou3J2a0VxFxKU06Y9PwzuHohO/SOS1ElV0fFKa2k5pBaOyDEhFpc8HkSj9qa5r9s
+510GolC5trZXMY+49dmH0QCHRxHqcLhMBJTS2Aq5JHT3SZsPxYo3MfTskAkFjId3WddpVh8+EnN
5Ksb1KrZ2TWQvle4/MZJeibL5tCq++MbLhfWpp/WZYct4pbmKd3mdyuzesQr8x3iQ/Bn+U5Fh0SO
gAVW/uoKauv8Q52ENZR0fCNHFzVxPIRyTP2cI40kQKCb+QMWEbXnMWtiH2wxh/WAn847v/XWNeUF
OTHWCiQkVoqjUdz/9dMuuWQRvPjawL/rWwKdmFaWsPuKgBhzV6RzanZ4DW8nu1PH6x5Hge0eh89r
VlW2vwxqL+cajfQLc9xloOQyQO4WeNI6el8/hBDByfpQsgUZjt/Nu3qztLDiAyBeqrTixcCdVJA8
4cm4IwgejtCnhxc2KUqfyvKRwOmT6uLS/9UEF1vz0Xn3wZkewUefnbE8MaSzWlWcCWSs1st84pJc
z9DwOE3OKKnaqa5vKCEfz5H6peAVCYgKzZC8VY+NRWKexbNZsCl1K5USsu6U0EU6Qas/+z4IYHu6
ZLD1vW0NWVj6MRsiFW3+EPA/
`protect end_protected
